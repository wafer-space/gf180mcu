VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__cor
  CLASS ENDCAP BOTTOMLEFT ;
  FOREIGN gf180mcu_fd_io__cor ;
  ORIGIN 0.000 0.000 ;
  SIZE 355.000 BY 355.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_COR_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 278.000 354.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 352.060 214.000 352.440 228.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.000 354.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.060 214.000 352.440 228.995 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 278.000 354.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 273.310 316.745 273.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 337.310 343.345 337.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.060 214.000 352.440 228.995 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.950 265.690 352.230 265.970 ;
      LAYER Metal5 ;
        RECT 351.950 265.690 352.230 265.970 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.910 270.000 352.290 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.920 278.000 352.300 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.945 294.000 352.325 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.010 334.000 352.390 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 214.000 350.740 229.000 351.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 265.310 313.415 265.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 281.310 320.060 281.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 297.310 326.710 297.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 209.310 289.930 209.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 188.320 283.200 188.700 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 118.000 350.800 125.000 351.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 140.320 263.145 140.700 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 156.320 269.835 156.700 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.040 350.980 172.320 351.260 ;
      LAYER Metal5 ;
        RECT 172.040 350.980 172.320 351.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.970 182.000 352.350 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.035 206.000 352.415 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 293.405 157.640 354.000 158.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.920 166.000 352.300 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.120 118.000 352.500 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 293.405 141.640 354.000 142.020 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 345.005 346.290 345.385 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 303.085 237.640 354.000 238.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.930 286.000 352.310 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.955 302.000 352.335 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.000 326.000 352.380 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.975 342.000 352.355 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 230.000 350.855 245.000 351.235 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 289.310 323.375 289.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 305.310 330.035 305.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 329.335 340.000 329.715 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 201.310 286.570 201.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 76.980 236.435 77.360 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 92.980 243.115 93.360 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 102.000 350.755 117.000 351.135 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 126.000 350.820 133.000 351.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 292.025 94.300 354.000 94.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.020 70.000 352.400 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.075 102.000 352.455 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 256.480 129.970 354.000 130.350 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.005 198.000 352.385 205.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.585 257.030 352.865 257.310 ;
      LAYER Metal5 ;
        RECT 352.585 257.030 352.865 257.310 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.965 310.000 352.345 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 257.310 310.075 257.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 313.310 333.350 313.690 354.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.580 249.690 352.860 249.970 ;
      LAYER Metal5 ;
        RECT 352.580 249.690 352.860 249.970 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.995 318.000 352.375 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 246.000 350.880 253.000 351.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 321.310 336.710 321.690 354.000 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 67.560 67.500 350.445 352.170 ;
      LAYER Metal1 ;
        RECT 65.540 65.540 355.000 355.000 ;
      LAYER Metal2 ;
        RECT 68.030 67.970 354.505 354.450 ;
      LAYER Metal3 ;
        RECT 85.300 353.700 85.700 354.450 ;
        RECT 101.300 353.700 101.700 354.450 ;
        RECT 117.300 353.700 117.700 354.450 ;
        RECT 125.300 353.700 125.700 354.450 ;
        RECT 133.300 353.700 133.700 354.450 ;
        RECT 149.300 353.700 149.700 354.450 ;
        RECT 165.300 353.700 165.700 354.450 ;
        RECT 181.300 353.700 181.700 354.450 ;
        RECT 197.300 353.700 197.700 354.450 ;
        RECT 205.300 353.700 205.700 354.450 ;
        RECT 213.300 353.700 213.700 354.450 ;
        RECT 229.300 353.700 229.700 354.450 ;
        RECT 245.300 353.700 245.700 354.450 ;
        RECT 253.300 353.700 253.700 354.450 ;
        RECT 261.300 353.700 261.700 354.450 ;
        RECT 269.300 353.700 269.700 354.450 ;
        RECT 277.300 353.700 277.700 354.450 ;
        RECT 285.300 353.700 285.700 354.450 ;
        RECT 293.300 353.700 293.700 354.450 ;
        RECT 301.300 353.700 301.700 354.450 ;
        RECT 309.300 353.700 309.700 354.450 ;
        RECT 317.300 353.700 317.700 354.450 ;
        RECT 325.300 353.700 325.700 354.450 ;
        RECT 333.300 353.700 333.700 354.450 ;
        RECT 341.300 353.700 341.700 354.450 ;
        RECT 348.690 353.700 355.000 354.450 ;
        RECT 70.000 348.690 355.000 353.700 ;
        RECT 70.000 341.700 353.700 348.690 ;
        RECT 70.000 341.300 355.000 341.700 ;
        RECT 70.000 333.700 353.700 341.300 ;
        RECT 70.000 333.300 355.000 333.700 ;
        RECT 70.000 325.700 353.700 333.300 ;
        RECT 70.000 325.300 355.000 325.700 ;
        RECT 70.000 317.700 353.700 325.300 ;
        RECT 70.000 317.300 355.000 317.700 ;
        RECT 70.000 309.700 353.700 317.300 ;
        RECT 70.000 309.300 355.000 309.700 ;
        RECT 70.000 301.700 353.700 309.300 ;
        RECT 70.000 301.300 355.000 301.700 ;
        RECT 70.000 293.700 353.700 301.300 ;
        RECT 70.000 293.300 355.000 293.700 ;
        RECT 70.000 285.700 353.700 293.300 ;
        RECT 70.000 285.300 355.000 285.700 ;
        RECT 70.000 277.700 353.700 285.300 ;
        RECT 70.000 277.300 355.000 277.700 ;
        RECT 70.000 269.700 353.700 277.300 ;
        RECT 70.000 269.300 355.000 269.700 ;
        RECT 70.000 261.700 353.700 269.300 ;
        RECT 70.000 261.300 355.000 261.700 ;
        RECT 70.000 253.700 353.700 261.300 ;
        RECT 70.000 253.300 355.000 253.700 ;
        RECT 70.000 245.700 353.700 253.300 ;
        RECT 70.000 245.300 355.000 245.700 ;
        RECT 70.000 229.700 353.700 245.300 ;
        RECT 70.000 229.295 355.000 229.700 ;
        RECT 70.000 213.700 351.760 229.295 ;
        RECT 352.740 213.700 355.000 229.295 ;
        RECT 70.000 213.300 355.000 213.700 ;
        RECT 70.000 205.700 353.700 213.300 ;
        RECT 70.000 205.300 355.000 205.700 ;
        RECT 70.000 197.700 353.700 205.300 ;
        RECT 70.000 197.300 355.000 197.700 ;
        RECT 70.000 181.700 353.700 197.300 ;
        RECT 70.000 181.300 355.000 181.700 ;
        RECT 70.000 165.700 353.700 181.300 ;
        RECT 70.000 165.300 355.000 165.700 ;
        RECT 70.000 149.700 353.700 165.300 ;
        RECT 70.000 149.300 355.000 149.700 ;
        RECT 70.000 133.700 353.700 149.300 ;
        RECT 70.000 133.300 355.000 133.700 ;
        RECT 70.000 125.700 353.700 133.300 ;
        RECT 70.000 125.300 355.000 125.700 ;
        RECT 70.000 117.700 353.700 125.300 ;
        RECT 70.000 117.300 355.000 117.700 ;
        RECT 70.000 101.700 353.700 117.300 ;
        RECT 70.000 101.300 355.000 101.700 ;
        RECT 70.000 85.700 353.700 101.300 ;
        RECT 70.000 85.300 355.000 85.700 ;
        RECT 70.000 70.000 353.700 85.300 ;
      LAYER Metal4 ;
        RECT 85.300 353.700 85.700 354.000 ;
        RECT 101.300 353.700 101.700 354.000 ;
        RECT 117.300 353.700 117.700 354.000 ;
        RECT 125.300 353.700 125.700 354.000 ;
        RECT 133.300 353.700 133.700 354.000 ;
        RECT 149.300 353.700 149.700 354.000 ;
        RECT 165.300 353.700 165.700 354.000 ;
        RECT 181.300 353.700 181.700 354.000 ;
        RECT 197.300 353.700 197.700 354.000 ;
        RECT 205.300 353.700 205.700 354.000 ;
        RECT 213.300 353.700 213.700 354.000 ;
        RECT 229.300 353.700 229.700 354.000 ;
        RECT 245.300 353.700 245.700 354.000 ;
        RECT 253.300 353.700 253.700 354.000 ;
        RECT 261.300 353.700 261.700 354.000 ;
        RECT 269.300 353.700 269.700 354.000 ;
        RECT 277.300 353.700 277.700 354.000 ;
        RECT 285.300 353.700 285.700 354.000 ;
        RECT 293.300 353.700 293.700 354.000 ;
        RECT 301.300 353.700 301.700 354.000 ;
        RECT 309.300 353.700 309.700 354.000 ;
        RECT 317.300 353.700 317.700 354.000 ;
        RECT 325.300 353.700 325.700 354.000 ;
        RECT 333.300 353.700 333.700 354.000 ;
        RECT 341.300 353.700 341.700 354.000 ;
        RECT 348.690 353.700 355.000 354.000 ;
        RECT 70.000 348.690 355.000 353.700 ;
        RECT 70.000 341.700 353.700 348.690 ;
        RECT 70.000 341.300 355.000 341.700 ;
        RECT 70.000 333.700 353.700 341.300 ;
        RECT 70.000 333.300 355.000 333.700 ;
        RECT 70.000 325.700 353.700 333.300 ;
        RECT 70.000 325.300 355.000 325.700 ;
        RECT 70.000 317.700 353.700 325.300 ;
        RECT 70.000 317.300 355.000 317.700 ;
        RECT 70.000 309.700 353.700 317.300 ;
        RECT 70.000 309.300 355.000 309.700 ;
        RECT 70.000 301.700 353.700 309.300 ;
        RECT 70.000 301.300 355.000 301.700 ;
        RECT 70.000 293.700 353.700 301.300 ;
        RECT 70.000 293.300 355.000 293.700 ;
        RECT 70.000 285.700 353.700 293.300 ;
        RECT 70.000 285.300 355.000 285.700 ;
        RECT 70.000 277.700 353.700 285.300 ;
        RECT 70.000 277.300 355.000 277.700 ;
        RECT 70.000 269.700 353.700 277.300 ;
        RECT 70.000 269.300 355.000 269.700 ;
        RECT 70.000 261.700 353.700 269.300 ;
        RECT 70.000 261.300 355.000 261.700 ;
        RECT 70.000 253.700 353.700 261.300 ;
        RECT 70.000 253.300 355.000 253.700 ;
        RECT 70.000 245.700 353.700 253.300 ;
        RECT 70.000 245.300 355.000 245.700 ;
        RECT 70.000 229.700 353.700 245.300 ;
        RECT 70.000 229.295 355.000 229.700 ;
        RECT 70.000 213.700 351.760 229.295 ;
        RECT 352.740 213.700 355.000 229.295 ;
        RECT 70.000 213.300 355.000 213.700 ;
        RECT 70.000 205.700 353.700 213.300 ;
        RECT 70.000 205.300 355.000 205.700 ;
        RECT 70.000 197.700 353.700 205.300 ;
        RECT 70.000 197.300 355.000 197.700 ;
        RECT 70.000 181.700 353.700 197.300 ;
        RECT 70.000 181.300 355.000 181.700 ;
        RECT 70.000 165.700 353.700 181.300 ;
        RECT 70.000 165.300 355.000 165.700 ;
        RECT 70.000 149.700 353.700 165.300 ;
        RECT 70.000 149.300 355.000 149.700 ;
        RECT 70.000 133.700 353.700 149.300 ;
        RECT 70.000 133.300 355.000 133.700 ;
        RECT 70.000 125.700 353.700 133.300 ;
        RECT 70.000 125.300 355.000 125.700 ;
        RECT 70.000 117.700 353.700 125.300 ;
        RECT 70.000 117.300 355.000 117.700 ;
        RECT 70.000 101.700 353.700 117.300 ;
        RECT 70.000 101.300 355.000 101.700 ;
        RECT 70.000 85.700 353.700 101.300 ;
        RECT 70.000 85.300 355.000 85.700 ;
        RECT 70.000 70.000 353.700 85.300 ;
      LAYER Metal5 ;
        RECT 348.890 353.500 355.000 354.000 ;
        RECT 70.000 235.935 76.480 353.500 ;
        RECT 77.860 242.615 92.480 353.500 ;
        RECT 93.860 351.700 139.820 353.500 ;
        RECT 93.860 351.680 125.500 351.700 ;
        RECT 93.860 351.635 117.500 351.680 ;
        RECT 93.860 350.255 101.500 351.635 ;
        RECT 133.500 350.320 139.820 351.700 ;
        RECT 125.500 350.300 139.820 350.320 ;
        RECT 117.500 350.255 139.820 350.300 ;
        RECT 93.860 262.645 139.820 350.255 ;
        RECT 141.200 269.335 155.820 353.500 ;
        RECT 157.200 351.760 187.820 353.500 ;
        RECT 157.200 350.480 171.540 351.760 ;
        RECT 172.820 350.480 187.820 351.760 ;
        RECT 157.200 282.700 187.820 350.480 ;
        RECT 189.200 286.070 200.810 353.500 ;
        RECT 202.190 289.430 208.810 353.500 ;
        RECT 210.190 351.760 256.810 353.500 ;
        RECT 210.190 351.735 245.500 351.760 ;
        RECT 210.190 351.620 229.500 351.735 ;
        RECT 210.190 350.240 213.500 351.620 ;
        RECT 253.500 350.380 256.810 351.760 ;
        RECT 245.500 350.355 256.810 350.380 ;
        RECT 229.500 350.240 256.810 350.355 ;
        RECT 210.190 309.575 256.810 350.240 ;
        RECT 258.190 312.915 264.810 353.500 ;
        RECT 266.190 316.245 272.810 353.500 ;
        RECT 274.190 319.560 280.810 353.500 ;
        RECT 282.190 322.875 288.810 353.500 ;
        RECT 290.190 326.210 296.810 353.500 ;
        RECT 298.190 329.535 304.810 353.500 ;
        RECT 306.190 332.850 312.810 353.500 ;
        RECT 314.190 336.210 320.810 353.500 ;
        RECT 322.190 339.500 328.835 353.500 ;
        RECT 330.215 342.845 336.810 353.500 ;
        RECT 338.190 345.790 344.505 353.500 ;
        RECT 345.885 348.890 355.000 353.500 ;
        RECT 345.885 345.790 351.475 348.890 ;
        RECT 338.190 342.845 351.475 345.790 ;
        RECT 330.215 341.500 351.475 342.845 ;
        RECT 352.855 341.500 353.500 348.890 ;
        RECT 330.215 339.500 351.510 341.500 ;
        RECT 322.190 336.210 351.510 339.500 ;
        RECT 314.190 333.500 351.510 336.210 ;
        RECT 352.890 333.500 353.500 341.500 ;
        RECT 314.190 332.850 351.500 333.500 ;
        RECT 306.190 329.535 351.500 332.850 ;
        RECT 298.190 326.210 351.500 329.535 ;
        RECT 290.190 325.500 351.500 326.210 ;
        RECT 352.880 325.500 353.500 333.500 ;
        RECT 290.190 322.875 351.495 325.500 ;
        RECT 282.190 319.560 351.495 322.875 ;
        RECT 274.190 317.500 351.495 319.560 ;
        RECT 352.875 317.500 353.500 325.500 ;
        RECT 274.190 316.245 351.465 317.500 ;
        RECT 266.190 312.915 351.465 316.245 ;
        RECT 258.190 309.575 351.465 312.915 ;
        RECT 210.190 309.500 351.465 309.575 ;
        RECT 352.845 309.500 353.500 317.500 ;
        RECT 210.190 301.500 351.455 309.500 ;
        RECT 352.835 301.500 353.500 309.500 ;
        RECT 210.190 293.500 351.445 301.500 ;
        RECT 352.825 293.500 353.500 301.500 ;
        RECT 210.190 289.430 351.430 293.500 ;
        RECT 202.190 286.070 351.430 289.430 ;
        RECT 189.200 285.500 351.430 286.070 ;
        RECT 352.810 285.500 353.500 293.500 ;
        RECT 189.200 282.700 351.420 285.500 ;
        RECT 157.200 277.500 351.420 282.700 ;
        RECT 352.800 277.500 353.500 285.500 ;
        RECT 157.200 269.500 351.410 277.500 ;
        RECT 352.790 269.500 353.500 277.500 ;
        RECT 157.200 269.335 353.500 269.500 ;
        RECT 141.200 266.470 353.500 269.335 ;
        RECT 141.200 265.190 351.450 266.470 ;
        RECT 352.730 265.190 353.500 266.470 ;
        RECT 141.200 262.645 353.500 265.190 ;
        RECT 93.860 257.810 353.500 262.645 ;
        RECT 93.860 256.530 352.085 257.810 ;
        RECT 353.365 256.530 353.500 257.810 ;
        RECT 93.860 250.470 353.500 256.530 ;
        RECT 93.860 249.190 352.080 250.470 ;
        RECT 353.360 249.190 353.500 250.470 ;
        RECT 93.860 242.615 353.500 249.190 ;
        RECT 77.860 238.520 353.500 242.615 ;
        RECT 77.860 237.140 302.585 238.520 ;
        RECT 77.860 235.935 353.500 237.140 ;
        RECT 70.000 229.500 353.500 235.935 ;
        RECT 70.000 229.495 355.000 229.500 ;
        RECT 70.000 213.500 351.560 229.495 ;
        RECT 352.940 213.500 355.000 229.495 ;
        RECT 70.000 205.500 351.535 213.500 ;
        RECT 352.915 205.500 353.500 213.500 ;
        RECT 70.000 197.500 351.505 205.500 ;
        RECT 352.885 197.500 353.500 205.500 ;
        RECT 70.000 181.500 351.470 197.500 ;
        RECT 352.850 181.500 353.500 197.500 ;
        RECT 70.000 165.500 351.420 181.500 ;
        RECT 352.800 165.500 353.500 181.500 ;
        RECT 70.000 158.520 353.500 165.500 ;
        RECT 70.000 157.140 292.905 158.520 ;
        RECT 70.000 142.520 353.500 157.140 ;
        RECT 70.000 141.140 292.905 142.520 ;
        RECT 70.000 130.850 353.500 141.140 ;
        RECT 70.000 129.470 255.980 130.850 ;
        RECT 70.000 125.500 353.500 129.470 ;
        RECT 70.000 117.500 351.620 125.500 ;
        RECT 353.000 117.500 353.500 125.500 ;
        RECT 70.000 101.500 351.575 117.500 ;
        RECT 352.955 101.500 353.500 117.500 ;
        RECT 70.000 95.180 353.500 101.500 ;
        RECT 70.000 93.800 291.525 95.180 ;
        RECT 70.000 85.500 353.500 93.800 ;
        RECT 70.000 70.000 351.520 85.500 ;
        RECT 352.900 70.000 353.500 85.500 ;
  END
END gf180mcu_fd_io__cor
END LIBRARY

