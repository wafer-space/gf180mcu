magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 758 870
<< pwell >>
rect -86 -86 758 352
<< metal1 >>
rect 0 724 672 844
rect 306 626 374 724
rect 141 326 318 438
rect 141 130 244 326
rect 497 320 591 676
rect 317 60 363 173
rect 466 115 591 320
rect 0 -60 672 60
<< obsm1 >>
rect 49 563 126 678
rect 49 516 451 563
rect 49 160 95 516
rect 394 366 451 516
<< labels >>
rlabel metal1 s 141 130 244 326 6 I
port 1 nsew default input
rlabel metal1 s 141 326 318 438 6 I
port 1 nsew default input
rlabel metal1 s 466 115 591 320 6 Z
port 2 nsew default output
rlabel metal1 s 497 320 591 676 6 Z
port 2 nsew default output
rlabel metal1 s 306 626 374 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 672 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 758 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 758 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 672 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 363 173 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1333148
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1330632
<< end >>
