magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -1030 29129 21660 29790
rect -1030 29053 21664 29129
rect -532 23867 21664 29053
rect -532 17407 21671 19961
<< mvpmos >>
rect -754 29194 -281 29649
rect -135 29194 338 29649
rect 484 29194 957 29649
rect 1103 29194 1576 29649
rect 1722 29194 2195 29649
rect 2341 29194 2814 29649
rect 2960 29194 3433 29649
rect 3579 29194 4052 29649
rect 4198 29194 4671 29649
rect 4817 29194 5290 29649
rect 5436 29194 5909 29649
rect 6055 29194 6528 29649
rect 6674 29194 7147 29649
rect 7293 29194 7766 29649
rect 7912 29194 8385 29649
rect 8531 29194 9004 29649
rect 9150 29194 9623 29649
rect 9769 29194 10242 29649
rect 10388 29194 10861 29649
rect 11007 29194 11480 29649
rect 11626 29194 12099 29649
rect 12245 29194 12718 29649
rect 12864 29194 13337 29649
rect 13483 29194 13956 29649
rect 14102 29194 14575 29649
rect 14721 29194 15194 29649
rect 15340 29194 15813 29649
rect 15959 29194 16432 29649
rect 16578 29194 17051 29649
rect 17197 29194 17670 29649
rect 17816 29194 18289 29649
rect 18435 29194 18908 29649
rect 19054 29194 19527 29649
rect 19673 29194 20146 29649
rect 20292 29194 20765 29649
rect 20911 29194 21384 29649
<< mvpdiff >>
rect -894 29604 -754 29649
rect -894 29558 -850 29604
rect -804 29558 -754 29604
rect -894 29286 -754 29558
rect -894 29240 -850 29286
rect -804 29240 -754 29286
rect -894 29194 -754 29240
rect -281 29604 -135 29649
rect -281 29558 -231 29604
rect -185 29558 -135 29604
rect -281 29286 -135 29558
rect -281 29240 -231 29286
rect -185 29240 -135 29286
rect -281 29194 -135 29240
rect 338 29604 484 29649
rect 338 29558 388 29604
rect 434 29558 484 29604
rect 338 29286 484 29558
rect 338 29240 388 29286
rect 434 29240 484 29286
rect 338 29194 484 29240
rect 957 29604 1103 29649
rect 957 29558 1007 29604
rect 1053 29558 1103 29604
rect 957 29286 1103 29558
rect 957 29240 1007 29286
rect 1053 29240 1103 29286
rect 957 29194 1103 29240
rect 1576 29604 1722 29649
rect 1576 29558 1626 29604
rect 1672 29558 1722 29604
rect 1576 29286 1722 29558
rect 1576 29240 1626 29286
rect 1672 29240 1722 29286
rect 1576 29194 1722 29240
rect 2195 29604 2341 29649
rect 2195 29558 2245 29604
rect 2291 29558 2341 29604
rect 2195 29286 2341 29558
rect 2195 29240 2245 29286
rect 2291 29240 2341 29286
rect 2195 29194 2341 29240
rect 2814 29604 2960 29649
rect 2814 29558 2864 29604
rect 2910 29558 2960 29604
rect 2814 29286 2960 29558
rect 2814 29240 2864 29286
rect 2910 29240 2960 29286
rect 2814 29194 2960 29240
rect 3433 29604 3579 29649
rect 3433 29558 3483 29604
rect 3529 29558 3579 29604
rect 3433 29286 3579 29558
rect 3433 29240 3483 29286
rect 3529 29240 3579 29286
rect 3433 29194 3579 29240
rect 4052 29604 4198 29649
rect 4052 29558 4102 29604
rect 4148 29558 4198 29604
rect 4052 29286 4198 29558
rect 4052 29240 4102 29286
rect 4148 29240 4198 29286
rect 4052 29194 4198 29240
rect 4671 29604 4817 29649
rect 4671 29558 4721 29604
rect 4767 29558 4817 29604
rect 4671 29286 4817 29558
rect 4671 29240 4721 29286
rect 4767 29240 4817 29286
rect 4671 29194 4817 29240
rect 5290 29604 5436 29649
rect 5290 29558 5340 29604
rect 5386 29558 5436 29604
rect 5290 29286 5436 29558
rect 5290 29240 5340 29286
rect 5386 29240 5436 29286
rect 5290 29194 5436 29240
rect 5909 29604 6055 29649
rect 5909 29558 5959 29604
rect 6005 29558 6055 29604
rect 5909 29286 6055 29558
rect 5909 29240 5959 29286
rect 6005 29240 6055 29286
rect 5909 29194 6055 29240
rect 6528 29604 6674 29649
rect 6528 29558 6578 29604
rect 6624 29558 6674 29604
rect 6528 29286 6674 29558
rect 6528 29240 6578 29286
rect 6624 29240 6674 29286
rect 6528 29194 6674 29240
rect 7147 29604 7293 29649
rect 7147 29558 7197 29604
rect 7243 29558 7293 29604
rect 7147 29286 7293 29558
rect 7147 29240 7197 29286
rect 7243 29240 7293 29286
rect 7147 29194 7293 29240
rect 7766 29604 7912 29649
rect 7766 29558 7816 29604
rect 7862 29558 7912 29604
rect 7766 29286 7912 29558
rect 7766 29240 7816 29286
rect 7862 29240 7912 29286
rect 7766 29194 7912 29240
rect 8385 29604 8531 29649
rect 8385 29558 8435 29604
rect 8481 29558 8531 29604
rect 8385 29286 8531 29558
rect 8385 29240 8435 29286
rect 8481 29240 8531 29286
rect 8385 29194 8531 29240
rect 9004 29604 9150 29649
rect 9004 29558 9054 29604
rect 9100 29558 9150 29604
rect 9004 29286 9150 29558
rect 9004 29240 9054 29286
rect 9100 29240 9150 29286
rect 9004 29194 9150 29240
rect 9623 29604 9769 29649
rect 9623 29558 9673 29604
rect 9719 29558 9769 29604
rect 9623 29286 9769 29558
rect 9623 29240 9673 29286
rect 9719 29240 9769 29286
rect 9623 29194 9769 29240
rect 10242 29604 10388 29649
rect 10242 29558 10292 29604
rect 10338 29558 10388 29604
rect 10242 29286 10388 29558
rect 10242 29240 10292 29286
rect 10338 29240 10388 29286
rect 10242 29194 10388 29240
rect 10861 29604 11007 29649
rect 10861 29558 10911 29604
rect 10957 29558 11007 29604
rect 10861 29286 11007 29558
rect 10861 29240 10911 29286
rect 10957 29240 11007 29286
rect 10861 29194 11007 29240
rect 11480 29604 11626 29649
rect 11480 29558 11530 29604
rect 11576 29558 11626 29604
rect 11480 29286 11626 29558
rect 11480 29240 11530 29286
rect 11576 29240 11626 29286
rect 11480 29194 11626 29240
rect 12099 29604 12245 29649
rect 12099 29558 12149 29604
rect 12195 29558 12245 29604
rect 12099 29286 12245 29558
rect 12099 29240 12149 29286
rect 12195 29240 12245 29286
rect 12099 29194 12245 29240
rect 12718 29604 12864 29649
rect 12718 29558 12768 29604
rect 12814 29558 12864 29604
rect 12718 29286 12864 29558
rect 12718 29240 12768 29286
rect 12814 29240 12864 29286
rect 12718 29194 12864 29240
rect 13337 29604 13483 29649
rect 13337 29558 13387 29604
rect 13433 29558 13483 29604
rect 13337 29286 13483 29558
rect 13337 29240 13387 29286
rect 13433 29240 13483 29286
rect 13337 29194 13483 29240
rect 13956 29604 14102 29649
rect 13956 29558 14006 29604
rect 14052 29558 14102 29604
rect 13956 29286 14102 29558
rect 13956 29240 14006 29286
rect 14052 29240 14102 29286
rect 13956 29194 14102 29240
rect 14575 29604 14721 29649
rect 14575 29558 14625 29604
rect 14671 29558 14721 29604
rect 14575 29286 14721 29558
rect 14575 29240 14625 29286
rect 14671 29240 14721 29286
rect 14575 29194 14721 29240
rect 15194 29604 15340 29649
rect 15194 29558 15244 29604
rect 15290 29558 15340 29604
rect 15194 29286 15340 29558
rect 15194 29240 15244 29286
rect 15290 29240 15340 29286
rect 15194 29194 15340 29240
rect 15813 29604 15959 29649
rect 15813 29558 15863 29604
rect 15909 29558 15959 29604
rect 15813 29286 15959 29558
rect 15813 29240 15863 29286
rect 15909 29240 15959 29286
rect 15813 29194 15959 29240
rect 16432 29604 16578 29649
rect 16432 29558 16482 29604
rect 16528 29558 16578 29604
rect 16432 29286 16578 29558
rect 16432 29240 16482 29286
rect 16528 29240 16578 29286
rect 16432 29194 16578 29240
rect 17051 29604 17197 29649
rect 17051 29558 17101 29604
rect 17147 29558 17197 29604
rect 17051 29286 17197 29558
rect 17051 29240 17101 29286
rect 17147 29240 17197 29286
rect 17051 29194 17197 29240
rect 17670 29604 17816 29649
rect 17670 29558 17720 29604
rect 17766 29558 17816 29604
rect 17670 29286 17816 29558
rect 17670 29240 17720 29286
rect 17766 29240 17816 29286
rect 17670 29194 17816 29240
rect 18289 29604 18435 29649
rect 18289 29558 18339 29604
rect 18385 29558 18435 29604
rect 18289 29286 18435 29558
rect 18289 29240 18339 29286
rect 18385 29240 18435 29286
rect 18289 29194 18435 29240
rect 18908 29604 19054 29649
rect 18908 29558 18958 29604
rect 19004 29558 19054 29604
rect 18908 29286 19054 29558
rect 18908 29240 18958 29286
rect 19004 29240 19054 29286
rect 18908 29194 19054 29240
rect 19527 29604 19673 29649
rect 19527 29558 19577 29604
rect 19623 29558 19673 29604
rect 19527 29286 19673 29558
rect 19527 29240 19577 29286
rect 19623 29240 19673 29286
rect 19527 29194 19673 29240
rect 20146 29604 20292 29649
rect 20146 29558 20196 29604
rect 20242 29558 20292 29604
rect 20146 29286 20292 29558
rect 20146 29240 20196 29286
rect 20242 29240 20292 29286
rect 20146 29194 20292 29240
rect 20765 29604 20911 29649
rect 20765 29558 20815 29604
rect 20861 29558 20911 29604
rect 20765 29286 20911 29558
rect 20765 29240 20815 29286
rect 20861 29240 20911 29286
rect 20765 29194 20911 29240
rect 21384 29604 21524 29649
rect 21384 29558 21434 29604
rect 21480 29558 21524 29604
rect 21384 29286 21524 29558
rect 21384 29240 21434 29286
rect 21480 29240 21524 29286
rect 21384 29194 21524 29240
<< mvpdiffc >>
rect -850 29558 -804 29604
rect -850 29240 -804 29286
rect -231 29558 -185 29604
rect -231 29240 -185 29286
rect 388 29558 434 29604
rect 388 29240 434 29286
rect 1007 29558 1053 29604
rect 1007 29240 1053 29286
rect 1626 29558 1672 29604
rect 1626 29240 1672 29286
rect 2245 29558 2291 29604
rect 2245 29240 2291 29286
rect 2864 29558 2910 29604
rect 2864 29240 2910 29286
rect 3483 29558 3529 29604
rect 3483 29240 3529 29286
rect 4102 29558 4148 29604
rect 4102 29240 4148 29286
rect 4721 29558 4767 29604
rect 4721 29240 4767 29286
rect 5340 29558 5386 29604
rect 5340 29240 5386 29286
rect 5959 29558 6005 29604
rect 5959 29240 6005 29286
rect 6578 29558 6624 29604
rect 6578 29240 6624 29286
rect 7197 29558 7243 29604
rect 7197 29240 7243 29286
rect 7816 29558 7862 29604
rect 7816 29240 7862 29286
rect 8435 29558 8481 29604
rect 8435 29240 8481 29286
rect 9054 29558 9100 29604
rect 9054 29240 9100 29286
rect 9673 29558 9719 29604
rect 9673 29240 9719 29286
rect 10292 29558 10338 29604
rect 10292 29240 10338 29286
rect 10911 29558 10957 29604
rect 10911 29240 10957 29286
rect 11530 29558 11576 29604
rect 11530 29240 11576 29286
rect 12149 29558 12195 29604
rect 12149 29240 12195 29286
rect 12768 29558 12814 29604
rect 12768 29240 12814 29286
rect 13387 29558 13433 29604
rect 13387 29240 13433 29286
rect 14006 29558 14052 29604
rect 14006 29240 14052 29286
rect 14625 29558 14671 29604
rect 14625 29240 14671 29286
rect 15244 29558 15290 29604
rect 15244 29240 15290 29286
rect 15863 29558 15909 29604
rect 15863 29240 15909 29286
rect 16482 29558 16528 29604
rect 16482 29240 16528 29286
rect 17101 29558 17147 29604
rect 17101 29240 17147 29286
rect 17720 29558 17766 29604
rect 17720 29240 17766 29286
rect 18339 29558 18385 29604
rect 18339 29240 18385 29286
rect 18958 29558 19004 29604
rect 18958 29240 19004 29286
rect 19577 29558 19623 29604
rect 19577 29240 19623 29286
rect 20196 29558 20242 29604
rect 20196 29240 20242 29286
rect 20815 29558 20861 29604
rect 20815 29240 20861 29286
rect 21434 29558 21480 29604
rect 21434 29240 21480 29286
<< polysilicon >>
rect -754 29803 -281 29858
rect -754 29757 -701 29803
rect -655 29757 -380 29803
rect -334 29757 -281 29803
rect -754 29649 -281 29757
rect -135 29803 338 29858
rect -135 29757 -82 29803
rect -36 29757 239 29803
rect 285 29757 338 29803
rect -135 29649 338 29757
rect 484 29803 957 29858
rect 484 29757 537 29803
rect 583 29757 858 29803
rect 904 29757 957 29803
rect 484 29649 957 29757
rect 1103 29803 1576 29858
rect 1103 29757 1156 29803
rect 1202 29757 1477 29803
rect 1523 29757 1576 29803
rect 1103 29649 1576 29757
rect 1722 29803 2195 29858
rect 1722 29757 1775 29803
rect 1821 29757 2096 29803
rect 2142 29757 2195 29803
rect 1722 29649 2195 29757
rect 2341 29803 2814 29858
rect 2341 29757 2394 29803
rect 2440 29757 2715 29803
rect 2761 29757 2814 29803
rect 2341 29649 2814 29757
rect 2960 29803 3433 29858
rect 2960 29757 3013 29803
rect 3059 29757 3334 29803
rect 3380 29757 3433 29803
rect 2960 29649 3433 29757
rect 3579 29803 4052 29858
rect 3579 29757 3632 29803
rect 3678 29757 3953 29803
rect 3999 29757 4052 29803
rect 3579 29649 4052 29757
rect 4198 29803 4671 29858
rect 4198 29757 4251 29803
rect 4297 29757 4572 29803
rect 4618 29757 4671 29803
rect 4198 29649 4671 29757
rect 4817 29803 5290 29858
rect 4817 29757 4870 29803
rect 4916 29757 5191 29803
rect 5237 29757 5290 29803
rect 4817 29649 5290 29757
rect 5436 29803 5909 29858
rect 5436 29757 5489 29803
rect 5535 29757 5810 29803
rect 5856 29757 5909 29803
rect 5436 29649 5909 29757
rect 6055 29803 6528 29858
rect 6055 29757 6108 29803
rect 6154 29757 6429 29803
rect 6475 29757 6528 29803
rect 6055 29649 6528 29757
rect 6674 29803 7147 29858
rect 6674 29757 6727 29803
rect 6773 29757 7048 29803
rect 7094 29757 7147 29803
rect 6674 29649 7147 29757
rect 7293 29803 7766 29858
rect 7293 29757 7346 29803
rect 7392 29757 7667 29803
rect 7713 29757 7766 29803
rect 7293 29649 7766 29757
rect 7912 29803 8385 29858
rect 7912 29757 7965 29803
rect 8011 29757 8286 29803
rect 8332 29757 8385 29803
rect 7912 29649 8385 29757
rect 8531 29803 9004 29858
rect 8531 29757 8584 29803
rect 8630 29757 8905 29803
rect 8951 29757 9004 29803
rect 8531 29649 9004 29757
rect 9150 29803 9623 29858
rect 9150 29757 9203 29803
rect 9249 29757 9524 29803
rect 9570 29757 9623 29803
rect 9150 29649 9623 29757
rect 9769 29803 10242 29858
rect 9769 29757 9822 29803
rect 9868 29757 10143 29803
rect 10189 29757 10242 29803
rect 9769 29649 10242 29757
rect 10388 29803 10861 29858
rect 10388 29757 10441 29803
rect 10487 29757 10762 29803
rect 10808 29757 10861 29803
rect 10388 29649 10861 29757
rect 11007 29803 11480 29858
rect 11007 29757 11060 29803
rect 11106 29757 11381 29803
rect 11427 29757 11480 29803
rect 11007 29649 11480 29757
rect 11626 29803 12099 29858
rect 11626 29757 11679 29803
rect 11725 29757 12000 29803
rect 12046 29757 12099 29803
rect 11626 29649 12099 29757
rect 12245 29803 12718 29858
rect 12245 29757 12298 29803
rect 12344 29757 12619 29803
rect 12665 29757 12718 29803
rect 12245 29649 12718 29757
rect 12864 29803 13337 29858
rect 12864 29757 12917 29803
rect 12963 29757 13238 29803
rect 13284 29757 13337 29803
rect 12864 29649 13337 29757
rect 13483 29803 13956 29858
rect 13483 29757 13536 29803
rect 13582 29757 13857 29803
rect 13903 29757 13956 29803
rect 13483 29649 13956 29757
rect 14102 29803 14575 29858
rect 14102 29757 14155 29803
rect 14201 29757 14476 29803
rect 14522 29757 14575 29803
rect 14102 29649 14575 29757
rect 14721 29803 15194 29858
rect 14721 29757 14774 29803
rect 14820 29757 15095 29803
rect 15141 29757 15194 29803
rect 14721 29649 15194 29757
rect 15340 29803 15813 29858
rect 15340 29757 15393 29803
rect 15439 29757 15714 29803
rect 15760 29757 15813 29803
rect 15340 29649 15813 29757
rect 15959 29803 16432 29858
rect 15959 29757 16012 29803
rect 16058 29757 16333 29803
rect 16379 29757 16432 29803
rect 15959 29649 16432 29757
rect 16578 29803 17051 29858
rect 16578 29757 16631 29803
rect 16677 29757 16952 29803
rect 16998 29757 17051 29803
rect 16578 29649 17051 29757
rect 17197 29803 17670 29858
rect 17197 29757 17250 29803
rect 17296 29757 17571 29803
rect 17617 29757 17670 29803
rect 17197 29649 17670 29757
rect 17816 29803 18289 29858
rect 17816 29757 17869 29803
rect 17915 29757 18190 29803
rect 18236 29757 18289 29803
rect 17816 29649 18289 29757
rect 18435 29803 18908 29858
rect 18435 29757 18488 29803
rect 18534 29757 18809 29803
rect 18855 29757 18908 29803
rect 18435 29649 18908 29757
rect 19054 29803 19527 29858
rect 19054 29757 19107 29803
rect 19153 29757 19428 29803
rect 19474 29757 19527 29803
rect 19054 29649 19527 29757
rect 19673 29803 20146 29858
rect 19673 29757 19726 29803
rect 19772 29757 20047 29803
rect 20093 29757 20146 29803
rect 19673 29649 20146 29757
rect 20292 29803 20765 29858
rect 20292 29757 20345 29803
rect 20391 29757 20666 29803
rect 20712 29757 20765 29803
rect 20292 29649 20765 29757
rect 20911 29803 21384 29858
rect 20911 29757 20964 29803
rect 21010 29757 21285 29803
rect 21331 29757 21384 29803
rect 20911 29649 21384 29757
rect -754 29112 -281 29194
rect -135 29112 338 29194
rect 484 29112 957 29194
rect 1103 29112 1576 29194
rect 1722 29112 2195 29194
rect 2341 29112 2814 29194
rect 2960 29112 3433 29194
rect 3579 29112 4052 29194
rect 4198 29112 4671 29194
rect 4817 29112 5290 29194
rect 5436 29112 5909 29194
rect 6055 29112 6528 29194
rect 6674 29112 7147 29194
rect 7293 29112 7766 29194
rect 7912 29112 8385 29194
rect 8531 29112 9004 29194
rect 9150 29112 9623 29194
rect 9769 29112 10242 29194
rect 10388 29112 10861 29194
rect 11007 29112 11480 29194
rect 11626 29112 12099 29194
rect 12245 29112 12718 29194
rect 12864 29112 13337 29194
rect 13483 29112 13956 29194
rect 14102 29112 14575 29194
rect 14721 29112 15194 29194
rect 15340 29112 15813 29194
rect 15959 29112 16432 29194
rect 16578 29112 17051 29194
rect 17197 29112 17670 29194
rect 17816 29112 18289 29194
rect 18435 29112 18908 29194
rect 19054 29112 19527 29194
rect 19673 29112 20146 29194
rect 20292 29112 20765 29194
rect 20911 29112 21384 29194
<< polycontact >>
rect -701 29757 -655 29803
rect -380 29757 -334 29803
rect -82 29757 -36 29803
rect 239 29757 285 29803
rect 537 29757 583 29803
rect 858 29757 904 29803
rect 1156 29757 1202 29803
rect 1477 29757 1523 29803
rect 1775 29757 1821 29803
rect 2096 29757 2142 29803
rect 2394 29757 2440 29803
rect 2715 29757 2761 29803
rect 3013 29757 3059 29803
rect 3334 29757 3380 29803
rect 3632 29757 3678 29803
rect 3953 29757 3999 29803
rect 4251 29757 4297 29803
rect 4572 29757 4618 29803
rect 4870 29757 4916 29803
rect 5191 29757 5237 29803
rect 5489 29757 5535 29803
rect 5810 29757 5856 29803
rect 6108 29757 6154 29803
rect 6429 29757 6475 29803
rect 6727 29757 6773 29803
rect 7048 29757 7094 29803
rect 7346 29757 7392 29803
rect 7667 29757 7713 29803
rect 7965 29757 8011 29803
rect 8286 29757 8332 29803
rect 8584 29757 8630 29803
rect 8905 29757 8951 29803
rect 9203 29757 9249 29803
rect 9524 29757 9570 29803
rect 9822 29757 9868 29803
rect 10143 29757 10189 29803
rect 10441 29757 10487 29803
rect 10762 29757 10808 29803
rect 11060 29757 11106 29803
rect 11381 29757 11427 29803
rect 11679 29757 11725 29803
rect 12000 29757 12046 29803
rect 12298 29757 12344 29803
rect 12619 29757 12665 29803
rect 12917 29757 12963 29803
rect 13238 29757 13284 29803
rect 13536 29757 13582 29803
rect 13857 29757 13903 29803
rect 14155 29757 14201 29803
rect 14476 29757 14522 29803
rect 14774 29757 14820 29803
rect 15095 29757 15141 29803
rect 15393 29757 15439 29803
rect 15714 29757 15760 29803
rect 16012 29757 16058 29803
rect 16333 29757 16379 29803
rect 16631 29757 16677 29803
rect 16952 29757 16998 29803
rect 17250 29757 17296 29803
rect 17571 29757 17617 29803
rect 17869 29757 17915 29803
rect 18190 29757 18236 29803
rect 18488 29757 18534 29803
rect 18809 29757 18855 29803
rect 19107 29757 19153 29803
rect 19428 29757 19474 29803
rect 19726 29757 19772 29803
rect 20047 29757 20093 29803
rect 20345 29757 20391 29803
rect 20666 29757 20712 29803
rect 20964 29757 21010 29803
rect 21285 29757 21331 29803
<< metal1 >>
rect -994 29890 -918 29900
rect -844 29890 -714 30180
rect 4539 29890 4703 30180
rect 9939 29900 10103 30180
rect 9791 29890 10103 29900
rect 15339 29890 15503 30180
rect 20739 29900 20903 30180
rect 20739 29890 21000 29900
rect -994 29888 21458 29890
rect -994 29732 -982 29888
rect -930 29803 9803 29888
rect 9959 29803 20832 29888
rect 20988 29803 21458 29888
rect -930 29757 -701 29803
rect -655 29757 -380 29803
rect -334 29757 -82 29803
rect -36 29757 239 29803
rect 285 29757 537 29803
rect 583 29757 858 29803
rect 904 29757 1156 29803
rect 1202 29757 1477 29803
rect 1523 29757 1775 29803
rect 1821 29757 2096 29803
rect 2142 29757 2394 29803
rect 2440 29757 2715 29803
rect 2761 29757 3013 29803
rect 3059 29757 3334 29803
rect 3380 29757 3632 29803
rect 3678 29757 3953 29803
rect 3999 29757 4251 29803
rect 4297 29757 4572 29803
rect 4618 29757 4870 29803
rect 4916 29757 5191 29803
rect 5237 29757 5489 29803
rect 5535 29757 5810 29803
rect 5856 29757 6108 29803
rect 6154 29757 6429 29803
rect 6475 29757 6727 29803
rect 6773 29757 7048 29803
rect 7094 29757 7346 29803
rect 7392 29757 7667 29803
rect 7713 29757 7965 29803
rect 8011 29757 8286 29803
rect 8332 29757 8584 29803
rect 8630 29757 8905 29803
rect 8951 29757 9203 29803
rect 9249 29757 9524 29803
rect 9570 29757 9803 29803
rect 9959 29757 10143 29803
rect 10189 29757 10441 29803
rect 10487 29757 10762 29803
rect 10808 29757 11060 29803
rect 11106 29757 11381 29803
rect 11427 29757 11679 29803
rect 11725 29757 12000 29803
rect 12046 29757 12298 29803
rect 12344 29757 12619 29803
rect 12665 29757 12917 29803
rect 12963 29757 13238 29803
rect 13284 29757 13536 29803
rect 13582 29757 13857 29803
rect 13903 29757 14155 29803
rect 14201 29757 14476 29803
rect 14522 29757 14774 29803
rect 14820 29757 15095 29803
rect 15141 29757 15393 29803
rect 15439 29757 15714 29803
rect 15760 29757 16012 29803
rect 16058 29757 16333 29803
rect 16379 29757 16631 29803
rect 16677 29757 16952 29803
rect 16998 29757 17250 29803
rect 17296 29757 17571 29803
rect 17617 29757 17869 29803
rect 17915 29757 18190 29803
rect 18236 29757 18488 29803
rect 18534 29757 18809 29803
rect 18855 29757 19107 29803
rect 19153 29757 19428 29803
rect 19474 29757 19726 29803
rect 19772 29757 20047 29803
rect 20093 29757 20345 29803
rect 20391 29757 20666 29803
rect 20712 29757 20832 29803
rect 21010 29757 21285 29803
rect 21331 29757 21458 29803
rect -930 29732 9803 29757
rect 9959 29732 20832 29757
rect 20988 29732 21458 29757
rect -994 29720 21458 29732
rect -885 29604 -769 29640
rect -885 29558 -850 29604
rect -804 29558 -769 29604
rect -885 29286 -769 29558
rect -885 29240 -850 29286
rect -804 29240 -769 29286
rect -885 28890 -769 29240
rect -266 29604 -150 29640
rect -266 29558 -231 29604
rect -185 29558 -150 29604
rect -266 29286 -150 29558
rect -266 29240 -231 29286
rect -185 29240 -150 29286
rect -266 28890 -150 29240
rect 353 29604 469 29640
rect 353 29558 388 29604
rect 434 29558 469 29604
rect 353 29286 469 29558
rect 353 29240 388 29286
rect 434 29240 469 29286
rect 353 28890 469 29240
rect 972 29604 1088 29640
rect 972 29558 1007 29604
rect 1053 29558 1088 29604
rect 972 29286 1088 29558
rect 972 29240 1007 29286
rect 1053 29240 1088 29286
rect 972 28890 1088 29240
rect 1591 29604 1707 29640
rect 1591 29558 1626 29604
rect 1672 29558 1707 29604
rect 1591 29286 1707 29558
rect 1591 29240 1626 29286
rect 1672 29240 1707 29286
rect 1591 28890 1707 29240
rect 2210 29604 2326 29640
rect 2210 29558 2245 29604
rect 2291 29558 2326 29604
rect 2210 29286 2326 29558
rect 2210 29240 2245 29286
rect 2291 29240 2326 29286
rect 2210 28890 2326 29240
rect 2829 29604 2945 29640
rect 2829 29558 2864 29604
rect 2910 29558 2945 29604
rect 2829 29286 2945 29558
rect 2829 29240 2864 29286
rect 2910 29240 2945 29286
rect 2829 28890 2945 29240
rect 3448 29604 3564 29640
rect 3448 29558 3483 29604
rect 3529 29558 3564 29604
rect 3448 29286 3564 29558
rect 3448 29240 3483 29286
rect 3529 29240 3564 29286
rect 3448 28890 3564 29240
rect 4067 29604 4183 29640
rect 4067 29558 4102 29604
rect 4148 29558 4183 29604
rect 4067 29286 4183 29558
rect 4067 29240 4102 29286
rect 4148 29240 4183 29286
rect 4067 28890 4183 29240
rect 4686 29604 4802 29640
rect 4686 29558 4721 29604
rect 4767 29558 4802 29604
rect 4686 29286 4802 29558
rect 4686 29240 4721 29286
rect 4767 29240 4802 29286
rect 4686 28890 4802 29240
rect 5305 29604 5421 29640
rect 5305 29558 5340 29604
rect 5386 29558 5421 29604
rect 5305 29286 5421 29558
rect 5305 29240 5340 29286
rect 5386 29240 5421 29286
rect 5305 28890 5421 29240
rect 5924 29604 6040 29640
rect 5924 29558 5959 29604
rect 6005 29558 6040 29604
rect 5924 29286 6040 29558
rect 5924 29240 5959 29286
rect 6005 29240 6040 29286
rect 5924 28890 6040 29240
rect 6543 29604 6659 29640
rect 6543 29558 6578 29604
rect 6624 29558 6659 29604
rect 6543 29286 6659 29558
rect 6543 29240 6578 29286
rect 6624 29240 6659 29286
rect 6543 28890 6659 29240
rect 7162 29604 7278 29640
rect 7162 29558 7197 29604
rect 7243 29558 7278 29604
rect 7162 29286 7278 29558
rect 7162 29240 7197 29286
rect 7243 29240 7278 29286
rect 7162 28890 7278 29240
rect 7781 29604 7897 29640
rect 7781 29558 7816 29604
rect 7862 29558 7897 29604
rect 7781 29286 7897 29558
rect 7781 29240 7816 29286
rect 7862 29240 7897 29286
rect 7781 28890 7897 29240
rect 8400 29604 8516 29640
rect 8400 29558 8435 29604
rect 8481 29558 8516 29604
rect 8400 29286 8516 29558
rect 8400 29240 8435 29286
rect 8481 29240 8516 29286
rect 8400 28890 8516 29240
rect 9019 29604 9135 29640
rect 9019 29558 9054 29604
rect 9100 29558 9135 29604
rect 9019 29286 9135 29558
rect 9019 29240 9054 29286
rect 9100 29240 9135 29286
rect 9019 28890 9135 29240
rect 9638 29604 9754 29640
rect 9638 29558 9673 29604
rect 9719 29558 9754 29604
rect 9638 29286 9754 29558
rect 9638 29240 9673 29286
rect 9719 29240 9754 29286
rect 9638 28890 9754 29240
rect 10257 29604 10373 29640
rect 10257 29558 10292 29604
rect 10338 29558 10373 29604
rect 10257 29286 10373 29558
rect 10257 29240 10292 29286
rect 10338 29240 10373 29286
rect 10257 28890 10373 29240
rect 10876 29604 10992 29640
rect 10876 29558 10911 29604
rect 10957 29558 10992 29604
rect 10876 29286 10992 29558
rect 10876 29240 10911 29286
rect 10957 29240 10992 29286
rect 10876 28890 10992 29240
rect 11495 29604 11611 29640
rect 11495 29558 11530 29604
rect 11576 29558 11611 29604
rect 11495 29286 11611 29558
rect 11495 29240 11530 29286
rect 11576 29240 11611 29286
rect 11495 28890 11611 29240
rect 12114 29604 12230 29640
rect 12114 29558 12149 29604
rect 12195 29558 12230 29604
rect 12114 29286 12230 29558
rect 12114 29240 12149 29286
rect 12195 29240 12230 29286
rect 12114 28890 12230 29240
rect 12733 29604 12849 29640
rect 12733 29558 12768 29604
rect 12814 29558 12849 29604
rect 12733 29286 12849 29558
rect 12733 29240 12768 29286
rect 12814 29240 12849 29286
rect 12733 28890 12849 29240
rect 13352 29604 13468 29640
rect 13352 29558 13387 29604
rect 13433 29558 13468 29604
rect 13352 29286 13468 29558
rect 13352 29240 13387 29286
rect 13433 29240 13468 29286
rect 13352 28890 13468 29240
rect 13971 29604 14087 29640
rect 13971 29558 14006 29604
rect 14052 29558 14087 29604
rect 13971 29286 14087 29558
rect 13971 29240 14006 29286
rect 14052 29240 14087 29286
rect 13971 28890 14087 29240
rect 14590 29604 14706 29640
rect 14590 29558 14625 29604
rect 14671 29558 14706 29604
rect 14590 29286 14706 29558
rect 14590 29240 14625 29286
rect 14671 29240 14706 29286
rect 14590 28890 14706 29240
rect 15209 29604 15325 29640
rect 15209 29558 15244 29604
rect 15290 29558 15325 29604
rect 15209 29286 15325 29558
rect 15209 29240 15244 29286
rect 15290 29240 15325 29286
rect 15209 28890 15325 29240
rect 15828 29604 15944 29640
rect 15828 29558 15863 29604
rect 15909 29558 15944 29604
rect 15828 29286 15944 29558
rect 15828 29240 15863 29286
rect 15909 29240 15944 29286
rect 15828 28890 15944 29240
rect 16447 29604 16563 29640
rect 16447 29558 16482 29604
rect 16528 29558 16563 29604
rect 16447 29286 16563 29558
rect 16447 29240 16482 29286
rect 16528 29240 16563 29286
rect 16447 28890 16563 29240
rect 17066 29604 17182 29640
rect 17066 29558 17101 29604
rect 17147 29558 17182 29604
rect 17066 29286 17182 29558
rect 17066 29240 17101 29286
rect 17147 29240 17182 29286
rect 17066 28890 17182 29240
rect 17685 29604 17801 29640
rect 17685 29558 17720 29604
rect 17766 29558 17801 29604
rect 17685 29286 17801 29558
rect 17685 29240 17720 29286
rect 17766 29240 17801 29286
rect 17685 28890 17801 29240
rect 18304 29604 18420 29640
rect 18304 29558 18339 29604
rect 18385 29558 18420 29604
rect 18304 29286 18420 29558
rect 18304 29240 18339 29286
rect 18385 29240 18420 29286
rect 18304 28890 18420 29240
rect 18923 29604 19039 29640
rect 18923 29558 18958 29604
rect 19004 29558 19039 29604
rect 18923 29286 19039 29558
rect 18923 29240 18958 29286
rect 19004 29240 19039 29286
rect 18923 28890 19039 29240
rect 19542 29604 19658 29640
rect 19542 29558 19577 29604
rect 19623 29558 19658 29604
rect 19542 29286 19658 29558
rect 19542 29240 19577 29286
rect 19623 29240 19658 29286
rect 19542 28890 19658 29240
rect 20161 29604 20277 29640
rect 20161 29558 20196 29604
rect 20242 29558 20277 29604
rect 20161 29286 20277 29558
rect 20161 29240 20196 29286
rect 20242 29240 20277 29286
rect 20161 28890 20277 29240
rect 20780 29604 20896 29640
rect 20780 29558 20815 29604
rect 20861 29558 20896 29604
rect 20780 29286 20896 29558
rect 20780 29240 20815 29286
rect 20861 29240 20896 29286
rect 20780 28890 20896 29240
rect 21399 29604 21515 29640
rect 21399 29558 21434 29604
rect 21480 29558 21515 29604
rect 21399 29286 21515 29558
rect 21399 29240 21434 29286
rect 21480 29240 21515 29286
rect 21399 28890 21515 29240
rect -885 28725 21515 28890
rect 14849 16092 15238 16230
rect 15664 16092 16243 16230
<< via1 >>
rect -982 29732 -930 29888
rect 9803 29803 9959 29888
rect 20832 29803 20988 29888
rect 9803 29757 9822 29803
rect 9822 29757 9868 29803
rect 9868 29757 9959 29803
rect 20832 29757 20964 29803
rect 20964 29757 20988 29803
rect 9803 29732 9959 29757
rect 20832 29732 20988 29757
<< metal2 >>
rect -1009 29987 -909 31176
rect -1009 29931 -983 29987
rect -927 29931 -909 29987
rect -1009 29888 -909 29931
rect -1009 29855 -982 29888
rect -930 29855 -909 29888
rect -1009 29799 -983 29855
rect -927 29799 -909 29855
rect -1009 29732 -982 29799
rect -930 29732 -909 29799
rect -1009 29723 -909 29732
rect -1009 29667 -983 29723
rect -927 29667 -909 29723
rect -1009 29591 -909 29667
rect -1009 29535 -983 29591
rect -927 29535 -909 29591
rect -1009 27521 -909 29535
rect -827 29107 -738 29955
rect -827 29069 -733 29107
rect -827 29013 -808 29069
rect -752 29013 -733 29069
rect -827 28883 -733 29013
rect -827 28827 -808 28883
rect -752 28827 -733 28883
rect -827 28788 -733 28827
rect -649 29072 -549 31176
rect -649 29016 -626 29072
rect -570 29016 -549 29072
rect -649 28940 -549 29016
rect -649 28884 -626 28940
rect -570 28884 -549 28940
rect -649 28808 -549 28884
rect -827 21746 -738 28788
rect -649 28752 -626 28808
rect -570 28752 -549 28808
rect -649 28676 -549 28752
rect -649 28620 -626 28676
rect -570 28620 -549 28676
rect -649 28544 -549 28620
rect -649 28488 -626 28544
rect -570 28488 -549 28544
rect -649 28412 -549 28488
rect -649 28356 -626 28412
rect -570 28356 -549 28412
rect -649 28280 -549 28356
rect -649 28224 -626 28280
rect -570 28224 -549 28280
rect -649 28148 -549 28224
rect -649 28092 -626 28148
rect -570 28092 -549 28148
rect -649 28016 -549 28092
rect -649 27960 -626 28016
rect -570 27960 -549 28016
rect -649 27884 -549 27960
rect -649 27828 -626 27884
rect -570 27828 -549 27884
rect -649 27752 -549 27828
rect -649 27696 -626 27752
rect -570 27696 -549 27752
rect -649 27620 -549 27696
rect -649 27564 -626 27620
rect -570 27564 -549 27620
rect -649 27516 -549 27564
rect 9791 29987 9891 31176
rect 9791 29931 9814 29987
rect 9870 29931 9891 29987
rect 9791 29900 9891 29931
rect 9791 29888 9971 29900
rect 9791 29732 9803 29888
rect 9959 29732 9971 29888
rect 9791 29723 9971 29732
rect 9791 29667 9814 29723
rect 9870 29720 9971 29723
rect 9870 29667 9891 29720
rect 9791 29591 9891 29667
rect 9791 29535 9814 29591
rect 9870 29535 9891 29591
rect 9791 27540 9891 29535
rect 10151 29072 10251 31176
rect 10151 29016 10177 29072
rect 10233 29016 10251 29072
rect 10151 28940 10251 29016
rect 10151 28884 10177 28940
rect 10233 28884 10251 28940
rect 10151 28808 10251 28884
rect 10151 28752 10177 28808
rect 10233 28752 10251 28808
rect 10151 28676 10251 28752
rect 10151 28620 10177 28676
rect 10233 28620 10251 28676
rect 10151 28544 10251 28620
rect 10151 28488 10177 28544
rect 10233 28488 10251 28544
rect 10151 28412 10251 28488
rect 10151 28356 10177 28412
rect 10233 28356 10251 28412
rect 10151 28280 10251 28356
rect 10151 28224 10177 28280
rect 10233 28224 10251 28280
rect 10151 28148 10251 28224
rect 10151 28092 10177 28148
rect 10233 28092 10251 28148
rect 10151 28016 10251 28092
rect 10151 27960 10177 28016
rect 10233 27960 10251 28016
rect 10151 27884 10251 27960
rect 10151 27828 10177 27884
rect 10233 27828 10251 27884
rect 10151 27752 10251 27828
rect 10151 27696 10177 27752
rect 10233 27696 10251 27752
rect 10151 27620 10251 27696
rect 10151 27564 10177 27620
rect 10233 27564 10251 27620
rect 10151 27539 10251 27564
rect 20591 29072 20691 31176
rect 20951 29987 21051 31176
rect 20951 29931 20975 29987
rect 21031 29931 21051 29987
rect 20951 29900 21051 29931
rect 20820 29888 21051 29900
rect 20820 29732 20832 29888
rect 20988 29855 21051 29888
rect 21031 29799 21051 29855
rect 20988 29732 21051 29799
rect 20820 29723 21051 29732
rect 20820 29720 20975 29723
rect 20591 29016 20612 29072
rect 20668 29016 20691 29072
rect 20591 28940 20691 29016
rect 20591 28884 20612 28940
rect 20668 28884 20691 28940
rect 20591 28808 20691 28884
rect 20591 28752 20612 28808
rect 20668 28752 20691 28808
rect 20591 28676 20691 28752
rect 20591 28620 20612 28676
rect 20668 28620 20691 28676
rect 20591 28544 20691 28620
rect 20591 28488 20612 28544
rect 20668 28488 20691 28544
rect 20591 28412 20691 28488
rect 20591 28356 20612 28412
rect 20668 28356 20691 28412
rect 20591 28280 20691 28356
rect 20591 28224 20612 28280
rect 20668 28224 20691 28280
rect 20591 28148 20691 28224
rect 20591 28092 20612 28148
rect 20668 28092 20691 28148
rect 20591 28016 20691 28092
rect 20591 27960 20612 28016
rect 20668 27960 20691 28016
rect 20591 27884 20691 27960
rect 20591 27828 20612 27884
rect 20668 27828 20691 27884
rect 20591 27752 20691 27828
rect 20591 27696 20612 27752
rect 20668 27696 20691 27752
rect 20591 27620 20691 27696
rect 20591 27564 20612 27620
rect 20668 27564 20691 27620
rect 20591 27524 20691 27564
rect 20951 29667 20975 29720
rect 21031 29667 21051 29723
rect 20951 29591 21051 29667
rect 20951 29535 20975 29591
rect 21031 29535 21051 29591
rect 20951 27527 21051 29535
<< via2 >>
rect -983 29931 -927 29987
rect -983 29799 -982 29855
rect -982 29799 -930 29855
rect -930 29799 -927 29855
rect -983 29667 -927 29723
rect -983 29535 -927 29591
rect -808 29013 -752 29069
rect -808 28827 -752 28883
rect -626 29016 -570 29072
rect -626 28884 -570 28940
rect -626 28752 -570 28808
rect -626 28620 -570 28676
rect -626 28488 -570 28544
rect -626 28356 -570 28412
rect -626 28224 -570 28280
rect -626 28092 -570 28148
rect -626 27960 -570 28016
rect -626 27828 -570 27884
rect -626 27696 -570 27752
rect -626 27564 -570 27620
rect 9814 29931 9870 29987
rect 9814 29799 9870 29855
rect 9814 29667 9870 29723
rect 9814 29535 9870 29591
rect 10177 29016 10233 29072
rect 10177 28884 10233 28940
rect 10177 28752 10233 28808
rect 10177 28620 10233 28676
rect 10177 28488 10233 28544
rect 10177 28356 10233 28412
rect 10177 28224 10233 28280
rect 10177 28092 10233 28148
rect 10177 27960 10233 28016
rect 10177 27828 10233 27884
rect 10177 27696 10233 27752
rect 10177 27564 10233 27620
rect 20975 29931 21031 29987
rect 20975 29799 20988 29855
rect 20988 29799 21031 29855
rect 20612 29016 20668 29072
rect 20612 28884 20668 28940
rect 20612 28752 20668 28808
rect 20612 28620 20668 28676
rect 20612 28488 20668 28544
rect 20612 28356 20668 28412
rect 20612 28224 20668 28280
rect 20612 28092 20668 28148
rect 20612 27960 20668 28016
rect 20612 27828 20668 27884
rect 20612 27696 20668 27752
rect 20612 27564 20668 27620
rect 20975 29667 21031 29723
rect 20975 29535 21031 29591
<< metal3 >>
rect -1115 38517 22810 38877
rect -1115 37737 22810 38097
rect -1115 36717 22810 37077
rect -1115 35937 22810 36297
rect -1115 34917 22810 35277
rect -1115 34137 22810 34497
rect -1115 33117 22810 33477
rect -1115 32337 22810 32697
rect -1115 31317 22810 31677
rect -1115 30537 22810 30897
rect -1186 29987 22164 29997
rect -1186 29931 -983 29987
rect -927 29931 9814 29987
rect 9870 29931 20975 29987
rect 21031 29931 22164 29987
rect -1186 29855 22164 29931
rect -1186 29799 -983 29855
rect -927 29799 9814 29855
rect 9870 29799 20975 29855
rect 21031 29799 22164 29855
rect -1186 29723 22164 29799
rect -1186 29667 -983 29723
rect -927 29667 9814 29723
rect 9870 29667 20975 29723
rect 21031 29667 22164 29723
rect -1186 29591 22164 29667
rect -1186 29535 -983 29591
rect -927 29535 9814 29591
rect 9870 29535 20975 29591
rect 21031 29535 22164 29591
rect -1186 29517 22164 29535
rect -826 29106 -733 29107
rect -1186 29072 22164 29106
rect -1186 29069 -626 29072
rect -1186 29013 -808 29069
rect -752 29016 -626 29069
rect -570 29016 10177 29072
rect 10233 29016 20612 29072
rect 20668 29016 22164 29072
rect -752 29013 22164 29016
rect -1186 28940 22164 29013
rect -1186 28884 -626 28940
rect -570 28884 10177 28940
rect 10233 28884 20612 28940
rect 20668 28884 22164 28940
rect -1186 28883 22164 28884
rect -1186 28827 -808 28883
rect -752 28827 22164 28883
rect -1186 28808 22164 28827
rect -1186 28752 -626 28808
rect -570 28752 10177 28808
rect 10233 28752 20612 28808
rect 20668 28752 22164 28808
rect -1186 28676 22164 28752
rect -1186 28620 -626 28676
rect -570 28620 10177 28676
rect 10233 28620 20612 28676
rect 20668 28620 22164 28676
rect -1186 28544 22164 28620
rect -1186 28488 -626 28544
rect -570 28488 10177 28544
rect 10233 28488 20612 28544
rect 20668 28488 22164 28544
rect -1186 28412 22164 28488
rect -1186 28356 -626 28412
rect -570 28356 10177 28412
rect 10233 28356 20612 28412
rect 20668 28356 22164 28412
rect -1186 28280 22164 28356
rect -1186 28224 -626 28280
rect -570 28224 10177 28280
rect 10233 28224 20612 28280
rect 20668 28224 22164 28280
rect -1186 28148 22164 28224
rect -1186 28092 -626 28148
rect -570 28092 10177 28148
rect 10233 28092 20612 28148
rect 20668 28092 22164 28148
rect -1186 28016 22164 28092
rect -1186 27960 -626 28016
rect -570 27960 10177 28016
rect 10233 27960 20612 28016
rect 20668 27960 22164 28016
rect -1186 27884 22164 27960
rect -1186 27828 -626 27884
rect -570 27828 10177 27884
rect 10233 27828 20612 27884
rect 20668 27828 22164 27884
rect -1186 27752 22164 27828
rect -1186 27696 -626 27752
rect -570 27696 10177 27752
rect 10233 27696 20612 27752
rect 20668 27696 22164 27752
rect -1186 27620 22164 27696
rect -1186 27564 -626 27620
rect -570 27564 10177 27620
rect 10233 27564 20612 27620
rect 20668 27564 22164 27620
rect -1186 27297 22164 27564
rect -672 21090 21329 21305
rect -672 20768 21329 20983
rect -672 20447 21329 20662
rect -672 20125 21329 20340
rect -672 19433 21329 19648
rect -672 19111 21329 19326
rect -672 18790 21329 19005
rect -672 18468 21329 18683
rect -672 17919 21329 18361
rect -672 16808 21329 17263
rect -672 12997 21329 15720
rect -672 11578 20757 12711
rect -672 9309 21329 11578
rect -701 8442 21329 9159
rect 20900 7827 21329 7828
rect -701 7017 21329 7827
rect -672 5155 21329 6472
rect -672 4929 20872 5005
rect -672 3134 21329 4496
rect -672 1961 21329 2576
rect -672 1285 21329 1854
rect -672 747 21329 1179
rect -672 155 21329 610
rect -709 -959 21420 -504
rect -709 -1598 21420 -1247
rect -709 -1810 21420 -1722
rect -709 -2041 21420 -1953
rect -709 -2517 21420 -2166
rect -709 -3242 21420 -2787
use col_64a_64x8m81_0  col_64a_64x8m81_0_0
timestamp 1755724134
transform 1 0 -1079 0 1 31107
box -68 -68 22268 7268
use dcap_103_novia_64x8m81  dcap_103_novia_64x8m81_0
array 0 35 619 0 0 0
timestamp 1755724134
transform 1 0 -827 0 1 29009
box 0 0 1 1
use ldummy_64x4_64x8m81  ldummy_64x4_64x8m81_0
timestamp 1755724134
transform 1 0 -541 0 1 30030
box -636 76 22573 9277
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_0
timestamp 1755724134
transform 1 0 -956 0 1 29810
box 0 0 1 1
use M2_M143105899832112_64x8m81  M2_M143105899832112_64x8m81_0
timestamp 1755724134
transform 1 0 9881 0 1 29810
box 0 0 1 1
use M2_M143105899832112_64x8m81  M2_M143105899832112_64x8m81_1
timestamp 1755724134
transform 1 0 20910 0 1 29810
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_0
timestamp 1755724134
transform 1 0 9842 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_1
timestamp 1755724134
transform 1 0 -955 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_2
timestamp 1755724134
transform 1 0 21003 0 1 29761
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_0
timestamp 1755724134
transform 1 0 20640 0 1 28318
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_1
timestamp 1755724134
transform 1 0 -598 0 1 28318
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_2
timestamp 1755724134
transform 1 0 10205 0 1 28318
box 0 0 1 1
use saout_m2_64x8m81  saout_m2_64x8m81_0
timestamp 1755724134
transform 1 0 -966 0 1 -1
box -269 -3393 7633 31140
use saout_m2_64x8m81  saout_m2_64x8m81_1
timestamp 1755724134
transform 1 0 9834 0 1 -1
box -269 -3393 7633 31140
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_0
timestamp 1755724134
transform -1 0 21008 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_1
timestamp 1755724134
transform -1 0 10208 0 1 6
box -269 -3400 7633 31133
use via2_x2_64x8m81  via2_x2_64x8m81_0
timestamp 1755724134
transform 1 0 -826 0 1 28789
box 0 0 1 1
<< labels >>
rlabel metal1 s 5690 15928 5690 15928 4 pcb[2]
port 1 nsew
rlabel metal1 s 3660 15928 3660 15928 4 pcb[3]
port 2 nsew
rlabel metal1 s 16496 15928 16496 15928 4 pcb[0]
port 3 nsew
rlabel metal1 s 14155 15928 14155 15928 4 pcb[1]
port 4 nsew
rlabel metal1 s 920 18163 920 18163 4 vdd
port 5 nsew
flabel metal1 s -808 31106 -808 31106 0 FreeSans 368 0 0 0 VDD
port 6 nsew
flabel metal1 s -367 -3355 -367 -3355 0 FreeSans 600 0 0 0 WEN[3]
port 7 nsew
flabel metal1 s 9597 -3329 9597 -3329 0 FreeSans 600 0 0 0 WEN[2]
port 8 nsew
flabel metal1 s 10395 -3329 10395 -3329 0 FreeSans 600 0 0 0 WEN[1]
port 9 nsew
flabel metal1 s 20398 -3329 20398 -3329 0 FreeSans 600 0 0 0 WEN[0]
port 10 nsew
rlabel metal1 s 16437 15928 16437 15928 4 pcb[0]
port 3 nsew
rlabel metal1 s 14224 15928 14224 15928 4 pcb[1]
port 4 nsew
rlabel metal1 s 3672 15928 3672 15928 4 pcb[3]
port 2 nsew
rlabel metal1 s 5615 15928 5615 15928 4 pcb[2]
port 1 nsew
flabel metal1 s -367 -3355 -367 -3355 0 FreeSans 600 0 0 0 WEN[3]
port 7 nsew
flabel metal1 s 9740 -3329 9740 -3329 0 FreeSans 600 0 0 0 WEN[2]
port 8 nsew
flabel metal1 s 10394 -3329 10394 -3329 0 FreeSans 600 0 0 0 WEN[1]
port 9 nsew
flabel metal1 s 20462 -3329 20462 -3329 0 FreeSans 600 0 0 0 WEN[0]
port 10 nsew
rlabel metal3 s 701 37868 701 37868 4 WL[7]
port 11 nsew
rlabel metal3 s 701 36968 701 36968 4 WL[6]
port 12 nsew
rlabel metal3 s 701 36068 701 36068 4 WL[5]
port 13 nsew
rlabel metal3 s 701 35168 701 35168 4 WL[4]
port 14 nsew
rlabel metal3 s 701 34268 701 34268 4 WL[3]
port 15 nsew
rlabel metal3 s 701 33368 701 33368 4 WL[2]
port 16 nsew
rlabel metal3 s 701 32468 701 32468 4 WL[1]
port 17 nsew
rlabel metal3 s 701 31568 701 31568 4 WL[0]
port 18 nsew
rlabel metal3 s 870 1467 870 1467 4 men
port 19 nsew
rlabel metal3 s 797 18592 797 18592 4 ypass[0]
port 20 nsew
rlabel metal3 s 797 18914 797 18914 4 ypass[1]
port 21 nsew
rlabel metal3 s 797 19231 797 19231 4 ypass[2]
port 22 nsew
rlabel metal3 s 797 19548 797 19548 4 ypass[3]
port 23 nsew
rlabel metal3 s 797 20204 797 20204 4 ypass[4]
port 24 nsew
rlabel metal3 s 797 20528 797 20528 4 ypass[5]
port 25 nsew
rlabel metal3 s 797 20845 797 20845 4 ypass[6]
port 26 nsew
rlabel metal3 s 797 21162 797 21162 4 ypass[7]
port 27 nsew
rlabel metal3 s 867 1467 867 1467 4 men
port 19 nsew
flabel metal3 s -334 8814 -334 8814 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 386 -334 386 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -305 1002 -305 1002 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 2322 -305 2322 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 5923 -305 5923 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 11468 -305 11468 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 22970 -305 22970 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 29782 -305 29782 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -334 3858 -334 3858 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 7580 -334 7580 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 14009 -334 14009 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 18141 -334 18141 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 27925 -334 27925 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 -708 -334 -708 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 -3027 -334 -3027 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -305 -1478 -305 -1478 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 -2341 -305 -2341 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s 793 -1999 793 -1999 0 FreeSans 448 0 0 0 GWEN
port 29 nsew
flabel metal3 s -325 4973 -325 4973 0 FreeSans 448 0 0 0 GWE
port 30 nsew
rlabel metal3 s -728 34270 -728 34270 4 WL[3]
port 15 nsew
rlabel metal3 s 797 18591 797 18591 4 ypass[0]
port 20 nsew
rlabel metal3 s 797 18913 797 18913 4 ypass[1]
port 21 nsew
rlabel metal3 s 797 19548 797 19548 4 ypass[3]
port 23 nsew
rlabel metal3 s 797 20203 797 20203 4 ypass[4]
port 24 nsew
rlabel metal3 s 797 20527 797 20527 4 ypass[5]
port 25 nsew
rlabel metal3 s 797 21162 797 21162 4 ypass[7]
port 27 nsew
rlabel metal3 s 868 1466 868 1466 4 men
port 19 nsew
flabel metal3 s -327 4977 -327 4977 0 FreeSans 448 0 0 0 GWE
port 30 nsew
flabel metal3 s -327 -3052 -327 -3052 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 -738 -327 -738 0 FreeSans 448 0 0 0 VDD
port 6 nsew
rlabel metal3 s -728 33370 -728 33370 4 WL[2]
port 16 nsew
rlabel metal3 s -728 32470 -728 32470 4 WL[1]
port 17 nsew
flabel metal3 s -327 390 -327 390 0 FreeSans 448 0 0 0 VDD
port 6 nsew
rlabel metal3 s -728 37870 -728 37870 4 WL[7]
port 11 nsew
rlabel metal3 s -728 36970 -728 36970 4 WL[6]
port 12 nsew
rlabel metal3 s -728 36070 -728 36070 4 WL[5]
port 13 nsew
rlabel metal3 s -728 35170 -728 35170 4 WL[4]
port 14 nsew
rlabel metal3 s -728 31570 -728 31570 4 WL[0]
port 18 nsew
rlabel metal3 s 798 20844 798 20844 4 ypass[6]
port 26 nsew
rlabel metal3 s 798 19230 798 19230 4 ypass[2]
port 22 nsew
flabel metal3 s -327 998 -327 998 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 2325 -327 2325 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 3859 -327 3859 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 7582 -327 7582 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 14010 -327 14010 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 18137 -327 18137 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 27926 -327 27926 0 FreeSans 448 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 29771 -327 29771 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 22970 -327 22970 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 11464 -327 11464 0 FreeSans 448 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 5924 -327 5924 0 FreeSans 448 0 0 0 VSS
port 28 nsew
rlabel metal2 s -454 104 -454 104 4 din[0]
port 31 nsew
rlabel metal2 s 9695 104 9695 104 4 din[1]
port 32 nsew
rlabel metal2 s 10331 104 10331 104 4 din[2]
port 33 nsew
rlabel metal2 s 8835 104 8835 104 4 q[1]
port 34 nsew
rlabel metal2 s 19234 29015 19234 29015 4 b[1]
port 35 nsew
rlabel metal2 s 17793 29015 17793 29015 4 b[4]
port 36 nsew
rlabel metal2 s 15518 29015 15518 29015 4 b[7]
port 37 nsew
rlabel metal2 s 14077 29015 14077 29015 4 b[10]
port 38 nsew
rlabel metal2 s 11802 29015 11802 29015 4 b[13]
port 39 nsew
rlabel metal2 s 9466 29015 9466 29015 4 b[16]
port 40 nsew
rlabel metal2 s 7190 29015 7190 29015 4 b[19]
port 41 nsew
rlabel metal2 s 5750 29015 5750 29015 4 b[22]
port 42 nsew
rlabel metal2 s 3475 29015 3475 29015 4 b[25]
port 43 nsew
rlabel metal2 s 2034 29015 2034 29015 4 b[28]
port 44 nsew
rlabel metal2 s -241 29015 -241 29015 4 b[31]
port 45 nsew
rlabel metal2 s 20495 104 20495 104 4 din[3]
port 46 nsew
rlabel metal2 s 382 104 382 104 4 q[0]
port 47 nsew
rlabel metal2 s 11187 104 11187 104 4 q[2]
port 48 nsew
rlabel metal2 s 19655 104 19655 104 4 q[3]
port 49 nsew
rlabel metal2 s 998 29015 998 29015 4 b[29]
port 50 nsew
rlabel metal2 s 3273 29015 3273 29015 4 b[26]
port 51 nsew
rlabel metal2 s 4713 29015 4713 29015 4 b[23]
port 52 nsew
rlabel metal2 s 6988 29015 6988 29015 4 b[20]
port 53 nsew
rlabel metal2 s 8429 29015 8429 29015 4 b[17]
port 54 nsew
rlabel metal2 s 11600 29015 11600 29015 4 b[14]
port 55 nsew
rlabel metal2 s 13041 29015 13041 29015 4 b[11]
port 56 nsew
rlabel metal2 s 15316 29015 15316 29015 4 b[8]
port 57 nsew
rlabel metal2 s 16757 29015 16757 29015 4 b[5]
port 58 nsew
rlabel metal2 s 19032 29015 19032 29015 4 b[2]
port 59 nsew
rlabel metal2 s 19853 29015 19853 29015 4 bb[0]
port 60 nsew
rlabel metal2 s 19651 29015 19651 29015 4 bb[1]
port 61 nsew
rlabel metal2 s 18614 29015 18614 29015 4 bb[2]
port 62 nsew
rlabel metal2 s 18412 29015 18412 29015 4 bb[3]
port 63 nsew
rlabel metal2 s 17376 29015 17376 29015 4 bb[4]
port 64 nsew
rlabel metal2 s 17174 29015 17174 29015 4 bb[5]
port 65 nsew
rlabel metal2 s 16137 29015 16137 29015 4 bb[6]
port 66 nsew
rlabel metal2 s 15935 29015 15935 29015 4 bb[7]
port 67 nsew
rlabel metal2 s 14899 29015 14899 29015 4 bb[8]
port 68 nsew
rlabel metal2 s 14697 29015 14697 29015 4 bb[9]
port 69 nsew
rlabel metal2 s 13660 29015 13660 29015 4 bb[10]
port 70 nsew
rlabel metal2 s 13458 29015 13458 29015 4 bb[11]
port 71 nsew
rlabel metal2 s 12422 29015 12422 29015 4 bb[12]
port 72 nsew
rlabel metal2 s 12220 29015 12220 29015 4 bb[13]
port 73 nsew
rlabel metal2 s 11183 29015 11183 29015 4 bb[14]
port 74 nsew
rlabel metal2 s 10981 29015 10981 29015 4 bb[15]
port 75 nsew
rlabel metal2 s 9048 29015 9048 29015 4 bb[16]
port 76 nsew
rlabel metal2 s 8846 29015 8846 29015 4 bb[17]
port 77 nsew
rlabel metal2 s 7810 29015 7810 29015 4 bb[18]
port 78 nsew
rlabel metal2 s 7608 29015 7608 29015 4 bb[19]
port 79 nsew
rlabel metal2 s 6571 29015 6571 29015 4 bb[20]
port 80 nsew
rlabel metal2 s 6369 29015 6369 29015 4 bb[21]
port 81 nsew
rlabel metal2 s 5333 29015 5333 29015 4 bb[22]
port 82 nsew
rlabel metal2 s 5131 29015 5131 29015 4 bb[23]
port 83 nsew
rlabel metal2 s 4094 29015 4094 29015 4 bb[24]
port 84 nsew
rlabel metal2 s 3892 29015 3892 29015 4 bb[25]
port 85 nsew
rlabel metal2 s 2856 29015 2856 29015 4 bb[26]
port 86 nsew
rlabel metal2 s 2654 29015 2654 29015 4 bb[27]
port 87 nsew
rlabel metal2 s 1617 29015 1617 29015 4 bb[28]
port 88 nsew
rlabel metal2 s 1415 29015 1415 29015 4 bb[29]
port 89 nsew
rlabel metal2 s 378 29015 378 29015 4 bb[30]
port 90 nsew
rlabel metal2 s 176 29015 176 29015 4 bb[31]
port 91 nsew
rlabel metal2 s 796 29015 796 29015 4 b[30]
port 92 nsew
rlabel metal2 s 2236 29015 2236 29015 4 b[27]
port 93 nsew
rlabel metal2 s 4511 29015 4511 29015 4 b[24]
port 94 nsew
rlabel metal2 s 10564 29015 10564 29015 4 b[15]
port 95 nsew
rlabel metal2 s 12839 29015 12839 29015 4 b[12]
port 96 nsew
rlabel metal2 s 14279 29015 14279 29015 4 b[9]
port 97 nsew
rlabel metal2 s 5952 29015 5952 29015 4 b[21]
port 98 nsew
rlabel metal2 s 20270 29015 20270 29015 4 b[0]
port 99 nsew
rlabel metal2 s 17995 29015 17995 29015 4 b[3]
port 100 nsew
rlabel metal2 s 16555 29015 16555 29015 4 b[6]
port 101 nsew
rlabel metal2 s 8227 29015 8227 29015 4 b[18]
port 102 nsew
rlabel metal3 701 38768 701 38768 4 WL[8]
rlabel metal3 -728 38770 -728 38770 4 WL[8]
<< properties >>
string FIXED_BBOX 15366 28635 15476 31202
string GDS_END 1646974
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1632750
string path 50.110 134.975 50.110 189.995 
<< end >>
