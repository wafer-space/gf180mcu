magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 3222 1094
<< pwell >>
rect -86 -86 3222 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 217 836 333
rect 884 217 1004 333
rect 1108 217 1228 333
rect 1276 217 1396 333
rect 1576 217 1696 333
rect 1800 217 1920 333
rect 2024 217 2144 333
rect 2192 217 2312 333
rect 2460 183 2580 333
rect 2828 69 2948 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 756 573 856 773
rect 904 573 1004 773
rect 1164 573 1264 773
rect 1312 573 1412 773
rect 1516 573 1616 773
rect 1720 573 1820 773
rect 2060 573 2160 773
rect 2212 573 2312 773
rect 2480 573 2580 793
rect 2828 573 2928 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 276 716 333
rect 628 230 641 276
rect 687 230 716 276
rect 628 217 716 230
rect 836 217 884 333
rect 1004 320 1108 333
rect 1004 274 1033 320
rect 1079 274 1108 320
rect 1004 217 1108 274
rect 1228 217 1276 333
rect 1396 217 1576 333
rect 1696 320 1800 333
rect 1696 274 1725 320
rect 1771 274 1800 320
rect 1696 217 1800 274
rect 1920 320 2024 333
rect 1920 274 1949 320
rect 1995 274 2024 320
rect 1920 217 2024 274
rect 2144 217 2192 333
rect 2312 242 2460 333
rect 2312 217 2385 242
rect 1456 127 1516 217
rect 1446 121 1516 127
rect 2372 196 2385 217
rect 2431 196 2460 242
rect 2372 183 2460 196
rect 2580 320 2668 333
rect 2580 274 2609 320
rect 2655 274 2668 320
rect 2580 183 2668 274
rect 2740 222 2828 333
rect 1446 114 1518 121
rect 1446 68 1459 114
rect 1505 68 1518 114
rect 2740 82 2753 222
rect 2799 82 2828 222
rect 2740 69 2828 82
rect 2948 320 3036 333
rect 2948 180 2977 320
rect 3023 180 3036 320
rect 2948 69 3036 180
rect 1446 55 1518 68
<< mvpdiff >>
rect 624 932 696 945
rect 56 836 144 849
rect 56 696 69 836
rect 115 696 144 836
rect 56 573 144 696
rect 244 836 348 849
rect 244 790 273 836
rect 319 790 348 836
rect 244 573 348 790
rect 448 632 536 849
rect 448 586 477 632
rect 523 586 536 632
rect 448 573 536 586
rect 624 792 637 932
rect 683 792 696 932
rect 2740 926 2828 939
rect 624 773 696 792
rect 2392 780 2480 793
rect 2392 773 2405 780
rect 624 573 756 773
rect 856 573 904 773
rect 1004 632 1164 773
rect 1004 586 1033 632
rect 1079 586 1164 632
rect 1004 573 1164 586
rect 1264 573 1312 773
rect 1412 760 1516 773
rect 1412 620 1441 760
rect 1487 620 1516 760
rect 1412 573 1516 620
rect 1616 726 1720 773
rect 1616 586 1645 726
rect 1691 586 1720 726
rect 1616 573 1720 586
rect 1820 726 2060 773
rect 1820 586 1949 726
rect 1995 586 2060 726
rect 1820 573 2060 586
rect 2160 573 2212 773
rect 2312 640 2405 773
rect 2451 640 2480 780
rect 2312 573 2480 640
rect 2580 726 2668 793
rect 2580 586 2609 726
rect 2655 586 2668 726
rect 2580 573 2668 586
rect 2740 786 2753 926
rect 2799 786 2828 926
rect 2740 573 2828 786
rect 2928 726 3016 939
rect 2928 586 2957 726
rect 3003 586 3016 726
rect 2928 573 3016 586
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 230 687 276
rect 1033 274 1079 320
rect 1725 274 1771 320
rect 1949 274 1995 320
rect 2385 196 2431 242
rect 2609 274 2655 320
rect 1459 68 1505 114
rect 2753 82 2799 222
rect 2977 180 3023 320
<< mvpdiffc >>
rect 69 696 115 836
rect 273 790 319 836
rect 477 586 523 632
rect 637 792 683 932
rect 1033 586 1079 632
rect 1441 620 1487 760
rect 1645 586 1691 726
rect 1949 586 1995 726
rect 2405 640 2451 780
rect 2609 586 2655 726
rect 2753 786 2799 926
rect 2957 586 3003 726
<< polysilicon >>
rect 2828 939 2928 983
rect 144 849 244 893
rect 348 849 448 893
rect 1164 865 1820 905
rect 1164 852 1264 865
rect 756 773 856 817
rect 904 773 1004 817
rect 1164 806 1177 852
rect 1223 806 1264 852
rect 1164 773 1264 806
rect 1312 773 1412 817
rect 1516 773 1616 817
rect 1720 773 1820 865
rect 2060 773 2160 817
rect 2212 773 2312 817
rect 2480 793 2580 837
rect 144 504 244 573
rect 144 458 157 504
rect 203 458 244 504
rect 144 377 244 458
rect 124 333 244 377
rect 348 433 448 573
rect 756 540 856 573
rect 756 494 769 540
rect 815 494 856 540
rect 756 481 856 494
rect 348 412 836 433
rect 348 366 361 412
rect 407 393 836 412
rect 407 366 468 393
rect 348 333 468 366
rect 716 333 836 393
rect 904 412 1004 573
rect 1164 529 1264 573
rect 904 377 926 412
rect 884 366 926 377
rect 972 366 1004 412
rect 1312 412 1412 573
rect 1516 540 1616 573
rect 1516 494 1529 540
rect 1575 494 1616 540
rect 1516 481 1616 494
rect 1312 393 1337 412
rect 884 333 1004 366
rect 1108 333 1228 377
rect 1276 366 1337 393
rect 1383 393 1412 412
rect 1383 366 1396 393
rect 1276 333 1396 366
rect 1576 377 1616 481
rect 1720 513 1820 573
rect 2060 540 2160 573
rect 2060 529 2101 540
rect 1720 473 2003 513
rect 2088 494 2101 529
rect 2147 494 2160 540
rect 2088 481 2160 494
rect 1963 439 2003 473
rect 1963 399 2064 439
rect 2024 377 2064 399
rect 2212 412 2312 573
rect 2212 377 2253 412
rect 1576 333 1696 377
rect 1800 333 1920 377
rect 2024 333 2144 377
rect 2192 366 2253 377
rect 2299 366 2312 412
rect 2480 540 2580 573
rect 2480 494 2493 540
rect 2539 494 2580 540
rect 2480 377 2580 494
rect 2192 333 2312 366
rect 2460 333 2580 377
rect 2828 412 2928 573
rect 2828 366 2841 412
rect 2887 377 2928 412
rect 2887 366 2948 377
rect 2828 333 2948 366
rect 124 131 244 175
rect 348 131 468 175
rect 716 173 836 217
rect 884 173 1004 217
rect 1108 184 1228 217
rect 1108 138 1121 184
rect 1167 138 1228 184
rect 1276 173 1396 217
rect 1108 125 1228 138
rect 1576 173 1696 217
rect 1800 184 1920 217
rect 1800 138 1813 184
rect 1859 138 1920 184
rect 2024 173 2144 217
rect 2192 173 2312 217
rect 2460 139 2580 183
rect 1800 125 1920 138
rect 2828 25 2948 69
<< polycontact >>
rect 1177 806 1223 852
rect 157 458 203 504
rect 769 494 815 540
rect 361 366 407 412
rect 926 366 972 412
rect 1529 494 1575 540
rect 1337 366 1383 412
rect 2101 494 2147 540
rect 2253 366 2299 412
rect 2493 494 2539 540
rect 2841 366 2887 412
rect 1121 138 1167 184
rect 1813 138 1859 184
<< metal1 >>
rect 0 932 3136 1098
rect 0 918 637 932
rect 69 836 115 847
rect 273 836 319 918
rect 273 779 319 790
rect 683 926 3136 932
rect 683 918 2753 926
rect 637 781 683 792
rect 1177 852 1223 863
rect 1177 735 1223 806
rect 388 731 1223 735
rect 115 696 1223 731
rect 69 689 1223 696
rect 1441 760 1487 918
rect 69 685 407 689
rect 142 504 315 542
rect 142 458 157 504
rect 203 458 315 504
rect 142 447 315 458
rect 361 412 407 685
rect 477 632 523 643
rect 477 551 523 586
rect 1033 632 1079 643
rect 2405 780 2451 918
rect 1441 609 1487 620
rect 1645 726 1691 737
rect 1033 551 1079 586
rect 477 540 815 551
rect 477 505 769 540
rect 49 366 361 401
rect 769 379 815 494
rect 1033 540 1575 551
rect 1033 494 1529 540
rect 1033 483 1575 494
rect 49 355 407 366
rect 49 320 95 355
rect 49 263 95 274
rect 497 333 815 379
rect 497 320 543 333
rect 497 263 543 274
rect 641 276 687 287
rect 273 234 319 245
rect 273 90 319 188
rect 641 90 687 230
rect 769 184 815 333
rect 926 412 978 423
rect 972 366 978 412
rect 926 242 978 366
rect 1033 320 1079 483
rect 1645 423 1691 586
rect 1337 412 1691 423
rect 1383 366 1691 412
rect 1337 355 1691 366
rect 1033 263 1079 274
rect 1645 331 1691 355
rect 1949 726 2359 737
rect 1995 691 2359 726
rect 1645 320 1771 331
rect 1645 274 1725 320
rect 1645 263 1771 274
rect 1949 320 1995 586
rect 1949 263 1995 274
rect 2101 540 2147 551
rect 2313 540 2359 691
rect 2799 918 3136 926
rect 2753 775 2799 786
rect 2405 629 2451 640
rect 2609 726 2655 737
rect 2313 494 2493 540
rect 2539 494 2550 540
rect 2101 217 2147 494
rect 2609 423 2655 586
rect 2942 726 3023 737
rect 2942 586 2957 726
rect 3003 586 3023 726
rect 2942 466 3023 586
rect 2253 412 2655 423
rect 2299 366 2841 412
rect 2887 366 2898 412
rect 2253 355 2655 366
rect 2609 320 2655 355
rect 2609 263 2655 274
rect 2977 320 3023 466
rect 1133 184 2147 217
rect 769 138 1121 184
rect 1167 171 1813 184
rect 1167 138 1178 171
rect 1802 138 1813 171
rect 1859 138 2147 184
rect 2385 242 2431 253
rect 1459 114 1505 125
rect 0 68 1459 90
rect 2385 90 2431 196
rect 2753 222 2799 233
rect 1505 82 2753 90
rect 2977 169 3023 180
rect 2799 82 3136 90
rect 1505 68 3136 82
rect 0 -90 3136 68
<< labels >>
flabel metal1 s 142 447 315 542 0 FreeSans 200 0 0 0 CLK
port 2 nsew clock input
flabel metal1 s 926 242 978 423 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 2942 466 3023 737 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3136 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 641 253 687 287 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 2977 169 3023 466 1 Q
port 3 nsew default output
rlabel metal1 s 2753 781 2799 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2405 781 2451 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1441 781 1487 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 637 781 683 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 781 319 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2753 779 2799 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2405 779 2451 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1441 779 1487 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 779 319 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2753 775 2799 779 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2405 775 2451 779 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1441 775 1487 779 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2405 629 2451 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1441 629 1487 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1441 609 1487 629 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2385 245 2431 253 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 245 687 253 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2385 233 2431 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2753 125 2799 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2385 125 2431 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 125 687 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2753 90 2799 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2385 90 2431 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1459 90 1505 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3136 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 1008
string GDS_END 587770
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 580324
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
