magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_0
timestamp 1755724134
transform 1 0 3990 0 1 9680
box 0 0 1 1
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_1
timestamp 1755724134
transform 1 0 6482 0 1 9680
box 0 0 1 1
use M1_PACTIVE_02_512x8m81  M1_PACTIVE_02_512x8m81_0
timestamp 1755724134
transform 1 0 5481 0 1 11376
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1755724134
transform 1 0 3314 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1755724134
transform 1 0 1522 0 1 3759
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1755724134
transform 1 0 2062 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1755724134
transform 1 0 3090 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_4
timestamp 1755724134
transform 1 0 494 0 1 3351
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_5
timestamp 1755724134
transform 1 0 1298 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_6
timestamp 1755724134
transform 1 0 270 0 1 3759
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_7
timestamp 1755724134
transform 1 0 2286 0 1 3351
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1755724134
transform 0 -1 4242 1 0 10079
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1755724134
transform 0 -1 5170 1 0 9970
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1755724134
transform 1 0 4928 0 1 10375
box 0 0 1 1
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1755724134
transform 1 0 5985 0 1 9417
box 0 0 1 1
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1755724134
transform 1 0 5455 0 1 9367
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1755724134
transform 1 0 7122 0 1 9979
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1755724134
transform 1 0 4267 0 1 9662
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1755724134
transform 1 0 6480 0 1 9676
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1755724134
transform 1 0 3991 0 1 9662
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1755724134
transform 1 0 4926 0 1 10469
box 0 0 1 1
use M2_M1$$43375660_R90_512x8m81  M2_M1$$43375660_R90_512x8m81_0
timestamp 1755724134
transform 0 -1 5457 1 0 9603
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1755724134
transform 1 0 4267 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1755724134
transform 1 0 4706 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1755724134
transform 1 0 6090 0 1 10519
box 0 0 1 1
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1755724134
transform 1 0 5169 0 1 3555
box 0 0 1 1
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_1
timestamp 1755724134
transform 1 0 6346 0 1 3353
box 0 0 1 1
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_2
timestamp 1755724134
transform 1 0 6860 0 1 3151
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1755724134
transform 1 0 4233 0 1 10076
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1755724134
transform 1 0 5161 0 1 10076
box 0 0 1 1
use M3_M2$$43368492_R90_512x8m81  M3_M2$$43368492_R90_512x8m81_0
timestamp 1755724134
transform 0 -1 5457 1 0 9603
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1755724134
transform 1 0 4267 0 1 9553
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1755724134
transform 1 0 6480 0 1 9567
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1755724134
transform 1 0 4267 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_3
timestamp 1755724134
transform 1 0 4706 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_4
timestamp 1755724134
transform 1 0 3991 0 1 9553
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_5
timestamp 1755724134
transform 1 0 6090 0 1 10519
box 0 0 1 1
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_0
timestamp 1755724134
transform 1 0 5951 0 1 10236
box -31 0 -30 1
use nmos_5p04310591302040_512x8m81  nmos_5p04310591302040_512x8m81_0
timestamp 1755724134
transform 1 0 4326 0 1 10240
box 0 0 1 1
use nmos_5p04310591302040_512x8m81  nmos_5p04310591302040_512x8m81_1
timestamp 1755724134
transform 1 0 4550 0 1 10240
box 0 0 1 1
use pmos_5p04310591302069_512x8m81  pmos_5p04310591302069_512x8m81_0
timestamp 1755724134
transform 1 0 5802 0 1 9519
box 0 0 1 1
use xpredec0_bot_512x8m81  xpredec0_bot_512x8m81_0
timestamp 1755724134
transform 1 0 5424 0 1 632
box -20 -633 1762 7949
use xpredec0_bot_512x8m81  xpredec0_bot_512x8m81_1
timestamp 1755724134
transform 1 0 3733 0 1 632
box -20 -633 1762 7949
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_0
timestamp 1755724134
transform -1 0 4025 0 1 34
box 441 438 1338 11038
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_1
timestamp 1755724134
transform -1 0 2233 0 1 34
box 441 438 1338 11038
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_2
timestamp 1755724134
transform 1 0 1351 0 1 34
box 441 438 1338 11038
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_3
timestamp 1755724134
transform 1 0 -441 0 1 34
box 441 438 1338 11038
<< properties >>
string GDS_END 957056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 949572
<< end >>
