magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 4342 870
<< pwell >>
rect -86 -86 4342 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2812 68 2932 232
rect 3036 68 3156 232
rect 3260 68 3380 232
rect 3484 68 3604 232
rect 3708 68 3828 232
rect 3932 68 4052 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
rect 3708 472 3808 716
rect 3932 472 4032 716
<< mvndiff >>
rect 36 142 124 232
rect 36 96 49 142
rect 95 96 124 142
rect 36 68 124 96
rect 244 192 348 232
rect 244 146 273 192
rect 319 146 348 192
rect 244 68 348 146
rect 468 142 572 232
rect 468 96 497 142
rect 543 96 572 142
rect 468 68 572 96
rect 692 192 796 232
rect 692 146 721 192
rect 767 146 796 192
rect 692 68 796 146
rect 916 142 1020 232
rect 916 96 945 142
rect 991 96 1020 142
rect 916 68 1020 96
rect 1140 192 1244 232
rect 1140 146 1169 192
rect 1215 146 1244 192
rect 1140 68 1244 146
rect 1364 142 1468 232
rect 1364 96 1393 142
rect 1439 96 1468 142
rect 1364 68 1468 96
rect 1588 192 1692 232
rect 1588 146 1617 192
rect 1663 146 1692 192
rect 1588 68 1692 146
rect 1812 142 1916 232
rect 1812 96 1841 142
rect 1887 96 1916 142
rect 1812 68 1916 96
rect 2036 192 2140 232
rect 2036 146 2065 192
rect 2111 146 2140 192
rect 2036 68 2140 146
rect 2260 142 2364 232
rect 2260 96 2289 142
rect 2335 96 2364 142
rect 2260 68 2364 96
rect 2484 192 2588 232
rect 2484 146 2513 192
rect 2559 146 2588 192
rect 2484 68 2588 146
rect 2708 142 2812 232
rect 2708 96 2737 142
rect 2783 96 2812 142
rect 2708 68 2812 96
rect 2932 192 3036 232
rect 2932 146 2961 192
rect 3007 146 3036 192
rect 2932 68 3036 146
rect 3156 142 3260 232
rect 3156 96 3185 142
rect 3231 96 3260 142
rect 3156 68 3260 96
rect 3380 192 3484 232
rect 3380 146 3409 192
rect 3455 146 3484 192
rect 3380 68 3484 146
rect 3604 142 3708 232
rect 3604 96 3633 142
rect 3679 96 3708 142
rect 3604 68 3708 96
rect 3828 192 3932 232
rect 3828 146 3857 192
rect 3903 146 3932 192
rect 3828 68 3932 146
rect 4052 142 4140 232
rect 4052 96 4081 142
rect 4127 96 4140 142
rect 4052 68 4140 96
<< mvpdiff >>
rect 36 665 124 716
rect 36 525 49 665
rect 95 525 124 665
rect 36 472 124 525
rect 224 665 348 716
rect 224 525 253 665
rect 299 525 348 665
rect 224 472 348 525
rect 448 665 572 716
rect 448 619 477 665
rect 523 619 572 665
rect 448 472 572 619
rect 672 665 796 716
rect 672 525 701 665
rect 747 525 796 665
rect 672 472 796 525
rect 896 665 1020 716
rect 896 619 925 665
rect 971 619 1020 665
rect 896 472 1020 619
rect 1120 665 1244 716
rect 1120 525 1149 665
rect 1195 525 1244 665
rect 1120 472 1244 525
rect 1344 665 1468 716
rect 1344 525 1373 665
rect 1419 525 1468 665
rect 1344 472 1468 525
rect 1568 665 1692 716
rect 1568 525 1617 665
rect 1663 525 1692 665
rect 1568 472 1692 525
rect 1792 691 1916 716
rect 1792 645 1821 691
rect 1867 645 1916 691
rect 1792 472 1916 645
rect 2016 665 2140 716
rect 2016 525 2045 665
rect 2091 525 2140 665
rect 2016 472 2140 525
rect 2240 691 2364 716
rect 2240 645 2269 691
rect 2315 645 2364 691
rect 2240 472 2364 645
rect 2464 665 2588 716
rect 2464 525 2493 665
rect 2539 525 2588 665
rect 2464 472 2588 525
rect 2688 691 2812 716
rect 2688 645 2717 691
rect 2763 645 2812 691
rect 2688 472 2812 645
rect 2912 665 3036 716
rect 2912 525 2941 665
rect 2987 525 3036 665
rect 2912 472 3036 525
rect 3136 691 3260 716
rect 3136 645 3165 691
rect 3211 645 3260 691
rect 3136 472 3260 645
rect 3360 665 3484 716
rect 3360 525 3389 665
rect 3435 525 3484 665
rect 3360 472 3484 525
rect 3584 691 3708 716
rect 3584 645 3613 691
rect 3659 645 3708 691
rect 3584 472 3708 645
rect 3808 665 3932 716
rect 3808 525 3837 665
rect 3883 525 3932 665
rect 3808 472 3932 525
rect 4032 665 4120 716
rect 4032 525 4061 665
rect 4107 525 4120 665
rect 4032 472 4120 525
<< mvndiffc >>
rect 49 96 95 142
rect 273 146 319 192
rect 497 96 543 142
rect 721 146 767 192
rect 945 96 991 142
rect 1169 146 1215 192
rect 1393 96 1439 142
rect 1617 146 1663 192
rect 1841 96 1887 142
rect 2065 146 2111 192
rect 2289 96 2335 142
rect 2513 146 2559 192
rect 2737 96 2783 142
rect 2961 146 3007 192
rect 3185 96 3231 142
rect 3409 146 3455 192
rect 3633 96 3679 142
rect 3857 146 3903 192
rect 4081 96 4127 142
<< mvpdiffc >>
rect 49 525 95 665
rect 253 525 299 665
rect 477 619 523 665
rect 701 525 747 665
rect 925 619 971 665
rect 1149 525 1195 665
rect 1373 525 1419 665
rect 1617 525 1663 665
rect 1821 645 1867 691
rect 2045 525 2091 665
rect 2269 645 2315 691
rect 2493 525 2539 665
rect 2717 645 2763 691
rect 2941 525 2987 665
rect 3165 645 3211 691
rect 3389 525 3435 665
rect 3613 645 3659 691
rect 3837 525 3883 665
rect 4061 525 4107 665
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 3708 716 3808 760
rect 3932 716 4032 760
rect 124 402 224 472
rect 348 402 448 472
rect 572 402 672 472
rect 796 402 896 472
rect 1020 402 1120 472
rect 1244 402 1344 472
rect 1468 407 1568 472
rect 1692 407 1792 472
rect 1916 407 2016 472
rect 2140 407 2240 472
rect 2364 407 2464 472
rect 2588 407 2688 472
rect 2812 407 2912 472
rect 3036 407 3136 472
rect 3260 407 3360 472
rect 3484 407 3584 472
rect 3708 407 3808 472
rect 3932 407 4032 472
rect 124 389 1364 402
rect 124 343 153 389
rect 1139 343 1364 389
rect 124 330 1364 343
rect 124 232 244 330
rect 348 232 468 330
rect 572 232 692 330
rect 796 232 916 330
rect 1020 300 1364 330
rect 1020 232 1140 300
rect 1244 232 1364 300
rect 1468 394 4052 407
rect 1468 348 1481 394
rect 2561 348 2925 394
rect 4005 348 4052 394
rect 1468 335 4052 348
rect 1468 232 1588 335
rect 1692 232 1812 335
rect 1916 232 2036 335
rect 2140 232 2260 335
rect 2364 232 2484 335
rect 2588 232 2708 335
rect 2812 232 2932 335
rect 3036 232 3156 335
rect 3260 232 3380 335
rect 3484 232 3604 335
rect 3708 232 3828 335
rect 3932 232 4052 335
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2812 24 2932 68
rect 3036 24 3156 68
rect 3260 24 3380 68
rect 3484 24 3604 68
rect 3708 24 3828 68
rect 3932 24 4052 68
<< polycontact >>
rect 153 343 1139 389
rect 1481 348 2561 394
rect 2925 348 4005 394
<< metal1 >>
rect 0 724 4256 844
rect 49 665 95 724
rect 49 506 95 525
rect 253 665 299 676
rect 477 665 523 724
rect 477 600 523 619
rect 701 665 747 676
rect 299 525 701 552
rect 925 665 971 724
rect 925 600 971 619
rect 1149 665 1195 676
rect 747 525 1149 552
rect 1373 665 1419 724
rect 1821 691 1867 724
rect 1195 525 1299 552
rect 253 506 1299 525
rect 1373 506 1419 525
rect 1617 665 1663 676
rect 2269 691 2315 724
rect 1821 634 1867 645
rect 2045 665 2091 676
rect 1663 525 2045 586
rect 2717 691 2763 724
rect 2269 634 2315 645
rect 2493 665 2539 676
rect 2091 525 2493 586
rect 3165 691 3211 724
rect 2717 634 2763 645
rect 2941 665 2987 676
rect 2539 525 2941 586
rect 3613 691 3659 724
rect 3165 634 3211 645
rect 3389 665 3435 676
rect 2987 525 3389 586
rect 3613 634 3659 645
rect 3837 665 3883 676
rect 3435 525 3837 586
rect 124 389 1140 430
rect 124 343 153 389
rect 1139 343 1140 389
rect 124 332 1140 343
rect 1252 405 1299 506
rect 1617 466 3883 525
rect 4061 665 4107 724
rect 4061 506 4107 525
rect 1252 394 2561 405
rect 1252 348 1481 394
rect 1252 337 2561 348
rect 1252 250 1299 337
rect 2664 284 2824 466
rect 2925 394 4052 406
rect 4005 348 4052 394
rect 2925 337 4052 348
rect 273 203 1299 250
rect 273 192 319 203
rect 38 142 106 153
rect 38 96 49 142
rect 95 96 106 142
rect 721 192 767 203
rect 273 135 319 146
rect 486 142 554 153
rect 38 60 106 96
rect 486 96 497 142
rect 543 96 554 142
rect 1169 192 1215 203
rect 721 135 767 146
rect 934 142 1002 153
rect 486 60 554 96
rect 934 96 945 142
rect 991 96 1002 142
rect 1617 196 3903 284
rect 1617 192 1669 196
rect 1169 135 1215 146
rect 1382 142 1450 153
rect 934 60 1002 96
rect 1382 96 1393 142
rect 1439 96 1450 142
rect 1663 146 1669 192
rect 1617 135 1669 146
rect 2065 192 2111 196
rect 1382 60 1450 96
rect 1830 96 1841 142
rect 1887 96 1898 142
rect 2065 135 2111 146
rect 2513 192 2559 196
rect 1830 60 1898 96
rect 2278 96 2289 142
rect 2335 96 2346 142
rect 2513 135 2559 146
rect 2961 192 3007 196
rect 2278 60 2346 96
rect 2726 96 2737 142
rect 2783 96 2794 142
rect 2961 135 3007 146
rect 3409 192 3455 196
rect 2726 60 2794 96
rect 3174 96 3185 142
rect 3231 96 3242 142
rect 3409 135 3455 146
rect 3857 192 3903 196
rect 3174 60 3242 96
rect 3622 96 3633 142
rect 3679 96 3690 142
rect 3857 106 3903 146
rect 4070 142 4138 153
rect 3622 60 3690 96
rect 4070 96 4081 142
rect 4127 96 4138 142
rect 4070 60 4138 96
rect 0 -60 4256 60
<< labels >>
flabel metal1 s 3837 586 3883 676 0 FreeSans 600 0 0 0 Z
port 2 nsew default output
flabel metal1 s 124 332 1140 430 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 4256 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 4070 142 4138 153 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 3389 586 3435 676 1 Z
port 2 nsew default output
rlabel metal1 s 2941 586 2987 676 1 Z
port 2 nsew default output
rlabel metal1 s 2493 586 2539 676 1 Z
port 2 nsew default output
rlabel metal1 s 2045 586 2091 676 1 Z
port 2 nsew default output
rlabel metal1 s 1617 586 1663 676 1 Z
port 2 nsew default output
rlabel metal1 s 1617 466 3883 586 1 Z
port 2 nsew default output
rlabel metal1 s 2664 284 2824 466 1 Z
port 2 nsew default output
rlabel metal1 s 1617 196 3903 284 1 Z
port 2 nsew default output
rlabel metal1 s 3857 135 3903 196 1 Z
port 2 nsew default output
rlabel metal1 s 3409 135 3455 196 1 Z
port 2 nsew default output
rlabel metal1 s 2961 135 3007 196 1 Z
port 2 nsew default output
rlabel metal1 s 2513 135 2559 196 1 Z
port 2 nsew default output
rlabel metal1 s 2065 135 2111 196 1 Z
port 2 nsew default output
rlabel metal1 s 1617 135 1669 196 1 Z
port 2 nsew default output
rlabel metal1 s 3857 106 3903 135 1 Z
port 2 nsew default output
rlabel metal1 s 4061 634 4107 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 634 3659 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 634 3211 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 634 2763 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 634 2315 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 634 1867 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 634 1419 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 634 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 634 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 634 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 600 4107 634 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 600 1419 634 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 600 971 634 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 600 523 634 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 600 95 634 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 506 4107 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 506 1419 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1382 142 1450 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 142 1002 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 142 554 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 142 106 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 142 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string GDS_END 1360632
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1351092
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
