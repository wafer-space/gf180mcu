magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
use via1_R90_512x8m81_0  via1_R90_512x8m81_0_0
timestamp 1755724134
transform 1 0 0 0 1 0
box 0 0 1 1
use via2_R90_512x8m81_0  via2_R90_512x8m81_0_0
timestamp 1755724134
transform 1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 612388
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 612296
<< end >>
