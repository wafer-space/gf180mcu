magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 7254 870
<< pwell >>
rect -86 -86 7254 352
<< mvnmos >>
rect 124 68 324 232
rect 572 68 772 232
rect 1020 68 1220 232
rect 1468 68 1668 232
rect 1916 68 2116 232
rect 2364 68 2564 232
rect 2812 68 3012 232
rect 3260 68 3460 232
rect 3708 68 3908 232
rect 4156 68 4356 232
rect 4604 68 4804 232
rect 5052 68 5252 232
rect 5500 68 5700 232
rect 5948 68 6148 232
rect 6396 68 6596 232
rect 6844 68 7044 232
<< mvpmos >>
rect 124 472 324 716
rect 572 472 772 716
rect 1020 472 1220 716
rect 1468 472 1668 716
rect 1916 472 2116 716
rect 2364 472 2564 716
rect 2812 472 3012 716
rect 3260 472 3460 716
rect 3708 472 3908 716
rect 4156 472 4356 716
rect 4604 472 4804 716
rect 5052 472 5252 716
rect 5500 472 5700 716
rect 5948 472 6148 716
rect 6396 472 6596 716
rect 6844 472 7044 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 324 192 412 232
rect 324 146 353 192
rect 399 146 412 192
rect 324 68 412 146
rect 484 192 572 232
rect 484 146 497 192
rect 543 146 572 192
rect 484 68 572 146
rect 772 192 860 232
rect 772 146 801 192
rect 847 146 860 192
rect 772 68 860 146
rect 932 192 1020 232
rect 932 146 945 192
rect 991 146 1020 192
rect 932 68 1020 146
rect 1220 192 1308 232
rect 1220 146 1249 192
rect 1295 146 1308 192
rect 1220 68 1308 146
rect 1380 192 1468 232
rect 1380 146 1393 192
rect 1439 146 1468 192
rect 1380 68 1468 146
rect 1668 192 1756 232
rect 1668 146 1697 192
rect 1743 146 1756 192
rect 1668 68 1756 146
rect 1828 192 1916 232
rect 1828 146 1841 192
rect 1887 146 1916 192
rect 1828 68 1916 146
rect 2116 192 2204 232
rect 2116 146 2145 192
rect 2191 146 2204 192
rect 2116 68 2204 146
rect 2276 192 2364 232
rect 2276 146 2289 192
rect 2335 146 2364 192
rect 2276 68 2364 146
rect 2564 192 2652 232
rect 2564 146 2593 192
rect 2639 146 2652 192
rect 2564 68 2652 146
rect 2724 192 2812 232
rect 2724 146 2737 192
rect 2783 146 2812 192
rect 2724 68 2812 146
rect 3012 192 3100 232
rect 3012 146 3041 192
rect 3087 146 3100 192
rect 3012 68 3100 146
rect 3172 192 3260 232
rect 3172 146 3185 192
rect 3231 146 3260 192
rect 3172 68 3260 146
rect 3460 192 3548 232
rect 3460 146 3489 192
rect 3535 146 3548 192
rect 3460 68 3548 146
rect 3620 192 3708 232
rect 3620 146 3633 192
rect 3679 146 3708 192
rect 3620 68 3708 146
rect 3908 192 3996 232
rect 3908 146 3937 192
rect 3983 146 3996 192
rect 3908 68 3996 146
rect 4068 192 4156 232
rect 4068 146 4081 192
rect 4127 146 4156 192
rect 4068 68 4156 146
rect 4356 192 4444 232
rect 4356 146 4385 192
rect 4431 146 4444 192
rect 4356 68 4444 146
rect 4516 192 4604 232
rect 4516 146 4529 192
rect 4575 146 4604 192
rect 4516 68 4604 146
rect 4804 192 4892 232
rect 4804 146 4833 192
rect 4879 146 4892 192
rect 4804 68 4892 146
rect 4964 192 5052 232
rect 4964 146 4977 192
rect 5023 146 5052 192
rect 4964 68 5052 146
rect 5252 192 5340 232
rect 5252 146 5281 192
rect 5327 146 5340 192
rect 5252 68 5340 146
rect 5412 192 5500 232
rect 5412 146 5425 192
rect 5471 146 5500 192
rect 5412 68 5500 146
rect 5700 192 5788 232
rect 5700 146 5729 192
rect 5775 146 5788 192
rect 5700 68 5788 146
rect 5860 192 5948 232
rect 5860 146 5873 192
rect 5919 146 5948 192
rect 5860 68 5948 146
rect 6148 192 6236 232
rect 6148 146 6177 192
rect 6223 146 6236 192
rect 6148 68 6236 146
rect 6308 192 6396 232
rect 6308 146 6321 192
rect 6367 146 6396 192
rect 6308 68 6396 146
rect 6596 192 6684 232
rect 6596 146 6625 192
rect 6671 146 6684 192
rect 6596 68 6684 146
rect 6756 192 6844 232
rect 6756 146 6769 192
rect 6815 146 6844 192
rect 6756 68 6844 146
rect 7044 192 7132 232
rect 7044 146 7073 192
rect 7119 146 7132 192
rect 7044 68 7132 146
<< mvpdiff >>
rect 36 657 124 716
rect 36 517 49 657
rect 95 517 124 657
rect 36 472 124 517
rect 324 657 412 716
rect 324 517 353 657
rect 399 517 412 657
rect 324 472 412 517
rect 484 657 572 716
rect 484 517 497 657
rect 543 517 572 657
rect 484 472 572 517
rect 772 657 860 716
rect 772 517 801 657
rect 847 517 860 657
rect 772 472 860 517
rect 932 657 1020 716
rect 932 517 945 657
rect 991 517 1020 657
rect 932 472 1020 517
rect 1220 657 1308 716
rect 1220 517 1249 657
rect 1295 517 1308 657
rect 1220 472 1308 517
rect 1380 657 1468 716
rect 1380 517 1393 657
rect 1439 517 1468 657
rect 1380 472 1468 517
rect 1668 657 1756 716
rect 1668 517 1697 657
rect 1743 517 1756 657
rect 1668 472 1756 517
rect 1828 657 1916 716
rect 1828 517 1841 657
rect 1887 517 1916 657
rect 1828 472 1916 517
rect 2116 657 2204 716
rect 2116 517 2145 657
rect 2191 517 2204 657
rect 2116 472 2204 517
rect 2276 657 2364 716
rect 2276 517 2289 657
rect 2335 517 2364 657
rect 2276 472 2364 517
rect 2564 657 2652 716
rect 2564 517 2593 657
rect 2639 517 2652 657
rect 2564 472 2652 517
rect 2724 657 2812 716
rect 2724 517 2737 657
rect 2783 517 2812 657
rect 2724 472 2812 517
rect 3012 657 3100 716
rect 3012 517 3041 657
rect 3087 517 3100 657
rect 3012 472 3100 517
rect 3172 657 3260 716
rect 3172 517 3185 657
rect 3231 517 3260 657
rect 3172 472 3260 517
rect 3460 657 3548 716
rect 3460 517 3489 657
rect 3535 517 3548 657
rect 3460 472 3548 517
rect 3620 657 3708 716
rect 3620 517 3633 657
rect 3679 517 3708 657
rect 3620 472 3708 517
rect 3908 657 3996 716
rect 3908 517 3937 657
rect 3983 517 3996 657
rect 3908 472 3996 517
rect 4068 657 4156 716
rect 4068 517 4081 657
rect 4127 517 4156 657
rect 4068 472 4156 517
rect 4356 657 4444 716
rect 4356 517 4385 657
rect 4431 517 4444 657
rect 4356 472 4444 517
rect 4516 657 4604 716
rect 4516 517 4529 657
rect 4575 517 4604 657
rect 4516 472 4604 517
rect 4804 657 4892 716
rect 4804 517 4833 657
rect 4879 517 4892 657
rect 4804 472 4892 517
rect 4964 657 5052 716
rect 4964 517 4977 657
rect 5023 517 5052 657
rect 4964 472 5052 517
rect 5252 657 5340 716
rect 5252 517 5281 657
rect 5327 517 5340 657
rect 5252 472 5340 517
rect 5412 657 5500 716
rect 5412 517 5425 657
rect 5471 517 5500 657
rect 5412 472 5500 517
rect 5700 657 5788 716
rect 5700 517 5729 657
rect 5775 517 5788 657
rect 5700 472 5788 517
rect 5860 657 5948 716
rect 5860 517 5873 657
rect 5919 517 5948 657
rect 5860 472 5948 517
rect 6148 657 6236 716
rect 6148 517 6177 657
rect 6223 517 6236 657
rect 6148 472 6236 517
rect 6308 657 6396 716
rect 6308 517 6321 657
rect 6367 517 6396 657
rect 6308 472 6396 517
rect 6596 657 6684 716
rect 6596 517 6625 657
rect 6671 517 6684 657
rect 6596 472 6684 517
rect 6756 657 6844 716
rect 6756 517 6769 657
rect 6815 517 6844 657
rect 6756 472 6844 517
rect 7044 657 7132 716
rect 7044 517 7073 657
rect 7119 517 7132 657
rect 7044 472 7132 517
<< mvndiffc >>
rect 49 146 95 192
rect 353 146 399 192
rect 497 146 543 192
rect 801 146 847 192
rect 945 146 991 192
rect 1249 146 1295 192
rect 1393 146 1439 192
rect 1697 146 1743 192
rect 1841 146 1887 192
rect 2145 146 2191 192
rect 2289 146 2335 192
rect 2593 146 2639 192
rect 2737 146 2783 192
rect 3041 146 3087 192
rect 3185 146 3231 192
rect 3489 146 3535 192
rect 3633 146 3679 192
rect 3937 146 3983 192
rect 4081 146 4127 192
rect 4385 146 4431 192
rect 4529 146 4575 192
rect 4833 146 4879 192
rect 4977 146 5023 192
rect 5281 146 5327 192
rect 5425 146 5471 192
rect 5729 146 5775 192
rect 5873 146 5919 192
rect 6177 146 6223 192
rect 6321 146 6367 192
rect 6625 146 6671 192
rect 6769 146 6815 192
rect 7073 146 7119 192
<< mvpdiffc >>
rect 49 517 95 657
rect 353 517 399 657
rect 497 517 543 657
rect 801 517 847 657
rect 945 517 991 657
rect 1249 517 1295 657
rect 1393 517 1439 657
rect 1697 517 1743 657
rect 1841 517 1887 657
rect 2145 517 2191 657
rect 2289 517 2335 657
rect 2593 517 2639 657
rect 2737 517 2783 657
rect 3041 517 3087 657
rect 3185 517 3231 657
rect 3489 517 3535 657
rect 3633 517 3679 657
rect 3937 517 3983 657
rect 4081 517 4127 657
rect 4385 517 4431 657
rect 4529 517 4575 657
rect 4833 517 4879 657
rect 4977 517 5023 657
rect 5281 517 5327 657
rect 5425 517 5471 657
rect 5729 517 5775 657
rect 5873 517 5919 657
rect 6177 517 6223 657
rect 6321 517 6367 657
rect 6625 517 6671 657
rect 6769 517 6815 657
rect 7073 517 7119 657
<< polysilicon >>
rect 124 716 324 760
rect 572 716 772 760
rect 1020 716 1220 760
rect 1468 716 1668 760
rect 1916 716 2116 760
rect 2364 716 2564 760
rect 2812 716 3012 760
rect 3260 716 3460 760
rect 3708 716 3908 760
rect 4156 716 4356 760
rect 4604 716 4804 760
rect 5052 716 5252 760
rect 5500 716 5700 760
rect 5948 716 6148 760
rect 6396 716 6596 760
rect 6844 716 7044 760
rect 124 438 324 472
rect 124 392 160 438
rect 300 392 324 438
rect 124 375 324 392
rect 572 438 772 472
rect 572 392 608 438
rect 748 392 772 438
rect 572 375 772 392
rect 1020 438 1220 472
rect 1020 392 1056 438
rect 1196 392 1220 438
rect 1020 375 1220 392
rect 1468 438 1668 472
rect 1468 392 1504 438
rect 1644 392 1668 438
rect 1468 375 1668 392
rect 1916 438 2116 472
rect 1916 392 1952 438
rect 2092 392 2116 438
rect 1916 375 2116 392
rect 2364 438 2564 472
rect 2364 392 2400 438
rect 2540 392 2564 438
rect 2364 375 2564 392
rect 2812 438 3012 472
rect 2812 392 2848 438
rect 2988 392 3012 438
rect 2812 375 3012 392
rect 3260 438 3460 472
rect 3260 392 3296 438
rect 3436 392 3460 438
rect 3260 375 3460 392
rect 3708 438 3908 472
rect 3708 392 3744 438
rect 3884 392 3908 438
rect 3708 375 3908 392
rect 4156 438 4356 472
rect 4156 392 4192 438
rect 4332 392 4356 438
rect 4156 375 4356 392
rect 4604 438 4804 472
rect 4604 392 4640 438
rect 4780 392 4804 438
rect 4604 375 4804 392
rect 5052 438 5252 472
rect 5052 392 5088 438
rect 5228 392 5252 438
rect 5052 375 5252 392
rect 5500 438 5700 472
rect 5500 392 5536 438
rect 5676 392 5700 438
rect 5500 375 5700 392
rect 5948 438 6148 472
rect 5948 392 5984 438
rect 6124 392 6148 438
rect 5948 375 6148 392
rect 6396 438 6596 472
rect 6396 392 6432 438
rect 6572 392 6596 438
rect 6396 375 6596 392
rect 6844 438 7044 472
rect 6844 392 6880 438
rect 7020 392 7044 438
rect 6844 375 7044 392
rect 124 311 324 324
rect 124 265 152 311
rect 292 265 324 311
rect 124 232 324 265
rect 572 311 772 324
rect 572 265 600 311
rect 740 265 772 311
rect 572 232 772 265
rect 1020 311 1220 324
rect 1020 265 1048 311
rect 1188 265 1220 311
rect 1020 232 1220 265
rect 1468 311 1668 324
rect 1468 265 1496 311
rect 1636 265 1668 311
rect 1468 232 1668 265
rect 1916 311 2116 324
rect 1916 265 1944 311
rect 2084 265 2116 311
rect 1916 232 2116 265
rect 2364 311 2564 324
rect 2364 265 2392 311
rect 2532 265 2564 311
rect 2364 232 2564 265
rect 2812 311 3012 324
rect 2812 265 2840 311
rect 2980 265 3012 311
rect 2812 232 3012 265
rect 3260 311 3460 324
rect 3260 265 3288 311
rect 3428 265 3460 311
rect 3260 232 3460 265
rect 3708 311 3908 324
rect 3708 265 3736 311
rect 3876 265 3908 311
rect 3708 232 3908 265
rect 4156 311 4356 324
rect 4156 265 4184 311
rect 4324 265 4356 311
rect 4156 232 4356 265
rect 4604 311 4804 324
rect 4604 265 4632 311
rect 4772 265 4804 311
rect 4604 232 4804 265
rect 5052 311 5252 324
rect 5052 265 5080 311
rect 5220 265 5252 311
rect 5052 232 5252 265
rect 5500 311 5700 324
rect 5500 265 5528 311
rect 5668 265 5700 311
rect 5500 232 5700 265
rect 5948 311 6148 324
rect 5948 265 5976 311
rect 6116 265 6148 311
rect 5948 232 6148 265
rect 6396 311 6596 324
rect 6396 265 6424 311
rect 6564 265 6596 311
rect 6396 232 6596 265
rect 6844 311 7044 324
rect 6844 265 6872 311
rect 7012 265 7044 311
rect 6844 232 7044 265
rect 124 24 324 68
rect 572 24 772 68
rect 1020 24 1220 68
rect 1468 24 1668 68
rect 1916 24 2116 68
rect 2364 24 2564 68
rect 2812 24 3012 68
rect 3260 24 3460 68
rect 3708 24 3908 68
rect 4156 24 4356 68
rect 4604 24 4804 68
rect 5052 24 5252 68
rect 5500 24 5700 68
rect 5948 24 6148 68
rect 6396 24 6596 68
rect 6844 24 7044 68
<< polycontact >>
rect 160 392 300 438
rect 608 392 748 438
rect 1056 392 1196 438
rect 1504 392 1644 438
rect 1952 392 2092 438
rect 2400 392 2540 438
rect 2848 392 2988 438
rect 3296 392 3436 438
rect 3744 392 3884 438
rect 4192 392 4332 438
rect 4640 392 4780 438
rect 5088 392 5228 438
rect 5536 392 5676 438
rect 5984 392 6124 438
rect 6432 392 6572 438
rect 6880 392 7020 438
rect 152 265 292 311
rect 600 265 740 311
rect 1048 265 1188 311
rect 1496 265 1636 311
rect 1944 265 2084 311
rect 2392 265 2532 311
rect 2840 265 2980 311
rect 3288 265 3428 311
rect 3736 265 3876 311
rect 4184 265 4324 311
rect 4632 265 4772 311
rect 5080 265 5220 311
rect 5528 265 5668 311
rect 5976 265 6116 311
rect 6424 265 6564 311
rect 6872 265 7012 311
<< metal1 >>
rect 0 724 7168 844
rect 49 657 95 678
rect 49 311 95 517
rect 353 657 399 724
rect 353 498 399 517
rect 497 657 543 678
rect 146 392 160 438
rect 300 392 399 438
rect 49 265 152 311
rect 292 265 304 311
rect 49 192 95 211
rect 49 60 95 146
rect 353 192 399 392
rect 497 311 543 517
rect 801 657 847 724
rect 801 498 847 517
rect 945 657 991 678
rect 594 392 608 438
rect 748 392 847 438
rect 497 265 600 311
rect 740 265 752 311
rect 353 106 399 146
rect 497 192 543 211
rect 497 60 543 146
rect 801 192 847 392
rect 945 311 991 517
rect 1249 657 1295 724
rect 1249 498 1295 517
rect 1393 657 1439 678
rect 1042 392 1056 438
rect 1196 392 1295 438
rect 945 265 1048 311
rect 1188 265 1200 311
rect 801 106 847 146
rect 945 192 991 211
rect 945 60 991 146
rect 1249 192 1295 392
rect 1393 311 1439 517
rect 1697 657 1743 724
rect 1697 498 1743 517
rect 1841 657 1887 678
rect 1490 392 1504 438
rect 1644 392 1743 438
rect 1393 265 1496 311
rect 1636 265 1648 311
rect 1249 106 1295 146
rect 1393 192 1439 211
rect 1393 60 1439 146
rect 1697 192 1743 392
rect 1841 311 1887 517
rect 2145 657 2191 724
rect 2145 498 2191 517
rect 2289 657 2335 678
rect 1938 392 1952 438
rect 2092 392 2191 438
rect 1841 265 1944 311
rect 2084 265 2096 311
rect 1697 106 1743 146
rect 1841 192 1887 211
rect 1841 60 1887 146
rect 2145 192 2191 392
rect 2289 311 2335 517
rect 2593 657 2639 724
rect 2593 498 2639 517
rect 2737 657 2783 678
rect 2386 392 2400 438
rect 2540 392 2639 438
rect 2289 265 2392 311
rect 2532 265 2544 311
rect 2145 106 2191 146
rect 2289 192 2335 211
rect 2289 60 2335 146
rect 2593 192 2639 392
rect 2737 311 2783 517
rect 3041 657 3087 724
rect 3041 498 3087 517
rect 3185 657 3231 678
rect 2834 392 2848 438
rect 2988 392 3087 438
rect 2737 265 2840 311
rect 2980 265 2992 311
rect 2593 106 2639 146
rect 2737 192 2783 211
rect 2737 60 2783 146
rect 3041 192 3087 392
rect 3185 311 3231 517
rect 3489 657 3535 724
rect 3489 498 3535 517
rect 3633 657 3679 678
rect 3282 392 3296 438
rect 3436 392 3535 438
rect 3185 265 3288 311
rect 3428 265 3440 311
rect 3041 106 3087 146
rect 3185 192 3231 211
rect 3185 60 3231 146
rect 3489 192 3535 392
rect 3633 311 3679 517
rect 3937 657 3983 724
rect 3937 498 3983 517
rect 4081 657 4127 678
rect 3730 392 3744 438
rect 3884 392 3983 438
rect 3633 265 3736 311
rect 3876 265 3888 311
rect 3489 106 3535 146
rect 3633 192 3679 211
rect 3633 60 3679 146
rect 3937 192 3983 392
rect 4081 311 4127 517
rect 4385 657 4431 724
rect 4385 498 4431 517
rect 4529 657 4575 678
rect 4178 392 4192 438
rect 4332 392 4431 438
rect 4081 265 4184 311
rect 4324 265 4336 311
rect 3937 106 3983 146
rect 4081 192 4127 211
rect 4081 60 4127 146
rect 4385 192 4431 392
rect 4529 311 4575 517
rect 4833 657 4879 724
rect 4833 498 4879 517
rect 4977 657 5023 678
rect 4626 392 4640 438
rect 4780 392 4879 438
rect 4529 265 4632 311
rect 4772 265 4784 311
rect 4385 106 4431 146
rect 4529 192 4575 211
rect 4529 60 4575 146
rect 4833 192 4879 392
rect 4977 311 5023 517
rect 5281 657 5327 724
rect 5281 498 5327 517
rect 5425 657 5471 678
rect 5074 392 5088 438
rect 5228 392 5327 438
rect 4977 265 5080 311
rect 5220 265 5232 311
rect 4833 106 4879 146
rect 4977 192 5023 211
rect 4977 60 5023 146
rect 5281 192 5327 392
rect 5425 311 5471 517
rect 5729 657 5775 724
rect 5729 498 5775 517
rect 5873 657 5919 678
rect 5522 392 5536 438
rect 5676 392 5775 438
rect 5425 265 5528 311
rect 5668 265 5680 311
rect 5281 106 5327 146
rect 5425 192 5471 211
rect 5425 60 5471 146
rect 5729 192 5775 392
rect 5873 311 5919 517
rect 6177 657 6223 724
rect 6177 498 6223 517
rect 6321 657 6367 678
rect 5970 392 5984 438
rect 6124 392 6223 438
rect 5873 265 5976 311
rect 6116 265 6128 311
rect 5729 106 5775 146
rect 5873 192 5919 211
rect 5873 60 5919 146
rect 6177 192 6223 392
rect 6321 311 6367 517
rect 6625 657 6671 724
rect 6625 498 6671 517
rect 6769 657 6815 678
rect 6418 392 6432 438
rect 6572 392 6671 438
rect 6321 265 6424 311
rect 6564 265 6576 311
rect 6177 106 6223 146
rect 6321 192 6367 211
rect 6321 60 6367 146
rect 6625 192 6671 392
rect 6769 311 6815 517
rect 7073 657 7119 724
rect 7073 498 7119 517
rect 6866 392 6880 438
rect 7020 392 7119 438
rect 6769 265 6872 311
rect 7012 265 7024 311
rect 6625 106 6671 146
rect 6769 192 6815 211
rect 6769 60 6815 146
rect 7073 192 7119 392
rect 7073 106 7119 146
rect 0 -60 7168 60
<< labels >>
flabel metal1 s 0 724 7168 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 6769 60 6815 211 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 7073 498 7119 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6625 498 6671 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6177 498 6223 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5729 498 5775 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5281 498 5327 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4833 498 4879 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4385 498 4431 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3937 498 3983 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3489 498 3535 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3041 498 3087 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2593 498 2639 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2145 498 2191 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 498 1743 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 498 1295 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 498 847 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6321 60 6367 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5873 60 5919 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5425 60 5471 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4977 60 5023 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 60 4575 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4081 60 4127 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3633 60 3679 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3185 60 3231 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2737 60 2783 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 211 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 7168 60 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 7168 784
string GDS_END 421994
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 402914
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
