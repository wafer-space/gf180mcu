magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 1318 1094
<< pwell >>
rect -86 -86 1318 453
<< metal1 >>
rect 0 918 1232 1098
rect 273 775 319 918
rect 27 451 203 542
rect 57 90 103 260
rect 251 242 418 413
rect 472 334 642 446
rect 690 433 866 542
rect 913 318 959 737
rect 1029 573 1208 654
rect 1029 483 1075 573
rect 913 288 1183 318
rect 485 242 1183 288
rect 485 215 531 242
rect 745 90 791 196
rect 1137 136 1183 242
rect 0 -90 1232 90
<< obsm1 >>
rect 709 826 1163 872
rect 69 634 115 750
rect 477 634 523 737
rect 709 710 755 826
rect 69 588 523 634
rect 477 575 523 588
rect 1117 710 1163 826
<< labels >>
rlabel metal1 s 1029 483 1075 573 6 A1
port 1 nsew default input
rlabel metal1 s 1029 573 1208 654 6 A1
port 1 nsew default input
rlabel metal1 s 690 433 866 542 6 A2
port 2 nsew default input
rlabel metal1 s 251 242 418 413 6 B1
port 3 nsew default input
rlabel metal1 s 27 451 203 542 6 B2
port 4 nsew default input
rlabel metal1 s 472 334 642 446 6 C
port 5 nsew default input
rlabel metal1 s 1137 136 1183 242 6 ZN
port 6 nsew default output
rlabel metal1 s 485 215 531 242 6 ZN
port 6 nsew default output
rlabel metal1 s 485 242 1183 288 6 ZN
port 6 nsew default output
rlabel metal1 s 913 288 1183 318 6 ZN
port 6 nsew default output
rlabel metal1 s 913 318 959 737 6 ZN
port 6 nsew default output
rlabel metal1 s 273 775 319 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 918 1232 1098 6 VDD
port 7 nsew power bidirectional abutment
rlabel nwell s -86 453 1318 1094 6 VNW
port 8 nsew power bidirectional
rlabel pwell s -86 -86 1318 453 6 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 0 -90 1232 90 8 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 745 90 791 196 6 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 57 90 103 260 6 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1232 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1219418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1215004
<< end >>
