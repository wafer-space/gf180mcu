magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< psubdiff >>
rect 70 96683 85816 96702
rect 70 96637 89 96683
rect 135 96637 213 96683
rect 259 96637 337 96683
rect 383 96637 461 96683
rect 507 96637 585 96683
rect 631 96637 709 96683
rect 755 96637 833 96683
rect 879 96637 957 96683
rect 1003 96637 1081 96683
rect 1127 96637 1205 96683
rect 1251 96637 1329 96683
rect 1375 96637 1453 96683
rect 1499 96637 1577 96683
rect 1623 96637 1701 96683
rect 1747 96637 1825 96683
rect 1871 96637 1949 96683
rect 1995 96637 2073 96683
rect 2119 96637 2197 96683
rect 2243 96637 2321 96683
rect 2367 96637 2445 96683
rect 2491 96637 2569 96683
rect 2615 96637 2693 96683
rect 2739 96637 2817 96683
rect 2863 96637 2941 96683
rect 2987 96637 3065 96683
rect 3111 96637 3189 96683
rect 3235 96637 3313 96683
rect 3359 96637 3437 96683
rect 3483 96637 3561 96683
rect 3607 96637 3685 96683
rect 3731 96637 3809 96683
rect 3855 96637 3933 96683
rect 3979 96637 4057 96683
rect 4103 96637 4181 96683
rect 4227 96637 4305 96683
rect 4351 96637 4429 96683
rect 4475 96637 4553 96683
rect 4599 96637 4677 96683
rect 4723 96637 4801 96683
rect 4847 96637 4925 96683
rect 4971 96637 5049 96683
rect 5095 96637 5173 96683
rect 5219 96637 5297 96683
rect 5343 96637 5421 96683
rect 5467 96637 5545 96683
rect 5591 96637 5669 96683
rect 5715 96637 5793 96683
rect 5839 96637 5917 96683
rect 5963 96637 6041 96683
rect 6087 96637 6165 96683
rect 6211 96637 6289 96683
rect 6335 96637 6413 96683
rect 6459 96637 6537 96683
rect 6583 96637 6661 96683
rect 6707 96637 6785 96683
rect 6831 96637 6909 96683
rect 6955 96637 7033 96683
rect 7079 96637 7157 96683
rect 7203 96637 7281 96683
rect 7327 96637 7405 96683
rect 7451 96637 7529 96683
rect 7575 96637 7653 96683
rect 7699 96637 7777 96683
rect 7823 96637 7901 96683
rect 7947 96637 8025 96683
rect 8071 96637 8149 96683
rect 8195 96637 8273 96683
rect 8319 96637 8397 96683
rect 8443 96637 8521 96683
rect 8567 96637 8645 96683
rect 8691 96637 8769 96683
rect 8815 96637 8893 96683
rect 8939 96637 9017 96683
rect 9063 96637 9141 96683
rect 9187 96637 9265 96683
rect 9311 96637 9389 96683
rect 9435 96637 9513 96683
rect 9559 96637 9637 96683
rect 9683 96637 9761 96683
rect 9807 96637 9885 96683
rect 9931 96637 10009 96683
rect 10055 96637 10133 96683
rect 10179 96637 10257 96683
rect 10303 96637 10381 96683
rect 10427 96637 10505 96683
rect 10551 96637 10629 96683
rect 10675 96637 10753 96683
rect 10799 96637 10877 96683
rect 10923 96637 11001 96683
rect 11047 96637 11125 96683
rect 11171 96637 11249 96683
rect 11295 96637 11373 96683
rect 11419 96637 11497 96683
rect 11543 96637 11621 96683
rect 11667 96637 11745 96683
rect 11791 96637 11869 96683
rect 11915 96637 11993 96683
rect 12039 96637 12117 96683
rect 12163 96637 12241 96683
rect 12287 96637 12365 96683
rect 12411 96637 12489 96683
rect 12535 96637 12613 96683
rect 12659 96637 12737 96683
rect 12783 96637 12861 96683
rect 12907 96637 12985 96683
rect 13031 96637 13109 96683
rect 13155 96637 13233 96683
rect 13279 96637 13357 96683
rect 13403 96637 13481 96683
rect 13527 96637 13605 96683
rect 13651 96637 13729 96683
rect 13775 96637 13853 96683
rect 13899 96637 13977 96683
rect 14023 96637 14101 96683
rect 14147 96637 14225 96683
rect 14271 96637 14349 96683
rect 14395 96637 14473 96683
rect 14519 96637 14597 96683
rect 14643 96637 14721 96683
rect 14767 96637 14845 96683
rect 14891 96637 14969 96683
rect 15015 96637 15093 96683
rect 15139 96637 15217 96683
rect 15263 96637 15341 96683
rect 15387 96637 15465 96683
rect 15511 96637 15589 96683
rect 15635 96637 15713 96683
rect 15759 96637 15837 96683
rect 15883 96637 15961 96683
rect 16007 96637 16085 96683
rect 16131 96637 16209 96683
rect 16255 96637 16333 96683
rect 16379 96637 16457 96683
rect 16503 96637 16581 96683
rect 16627 96637 16705 96683
rect 16751 96637 16829 96683
rect 16875 96637 16953 96683
rect 16999 96637 17077 96683
rect 17123 96637 17201 96683
rect 17247 96637 17325 96683
rect 17371 96637 17449 96683
rect 17495 96637 17573 96683
rect 17619 96637 17697 96683
rect 17743 96637 17821 96683
rect 17867 96637 17945 96683
rect 17991 96637 18069 96683
rect 18115 96637 18193 96683
rect 18239 96637 18317 96683
rect 18363 96637 18441 96683
rect 18487 96637 18565 96683
rect 18611 96637 18689 96683
rect 18735 96637 18813 96683
rect 18859 96637 18937 96683
rect 18983 96637 19061 96683
rect 19107 96637 19185 96683
rect 19231 96637 19309 96683
rect 19355 96637 19433 96683
rect 19479 96637 19557 96683
rect 19603 96637 19681 96683
rect 19727 96637 19805 96683
rect 19851 96637 19929 96683
rect 19975 96637 20053 96683
rect 20099 96637 20177 96683
rect 20223 96637 20301 96683
rect 20347 96637 20425 96683
rect 20471 96637 20549 96683
rect 20595 96637 20673 96683
rect 20719 96637 20797 96683
rect 20843 96637 20921 96683
rect 20967 96637 21045 96683
rect 21091 96637 21169 96683
rect 21215 96637 21293 96683
rect 21339 96637 21417 96683
rect 21463 96637 21541 96683
rect 21587 96637 21665 96683
rect 21711 96637 21789 96683
rect 21835 96637 21913 96683
rect 21959 96637 22037 96683
rect 22083 96637 22161 96683
rect 22207 96637 22285 96683
rect 22331 96637 22409 96683
rect 22455 96637 22533 96683
rect 22579 96637 22657 96683
rect 22703 96637 22781 96683
rect 22827 96637 22905 96683
rect 22951 96637 23029 96683
rect 23075 96637 23153 96683
rect 23199 96637 23277 96683
rect 23323 96637 23401 96683
rect 23447 96637 23525 96683
rect 23571 96637 23649 96683
rect 23695 96637 23773 96683
rect 23819 96637 23897 96683
rect 23943 96637 24021 96683
rect 24067 96637 24145 96683
rect 24191 96637 24269 96683
rect 24315 96637 24393 96683
rect 24439 96637 24517 96683
rect 24563 96637 24641 96683
rect 24687 96637 24765 96683
rect 24811 96637 24889 96683
rect 24935 96637 25013 96683
rect 25059 96637 25137 96683
rect 25183 96637 25261 96683
rect 25307 96637 25385 96683
rect 25431 96637 25509 96683
rect 25555 96637 25633 96683
rect 25679 96637 25757 96683
rect 25803 96637 25881 96683
rect 25927 96637 26005 96683
rect 26051 96637 26129 96683
rect 26175 96637 26253 96683
rect 26299 96637 26377 96683
rect 26423 96637 26501 96683
rect 26547 96637 26625 96683
rect 26671 96637 26749 96683
rect 26795 96637 26873 96683
rect 26919 96637 26997 96683
rect 27043 96637 27121 96683
rect 27167 96637 27245 96683
rect 27291 96637 27369 96683
rect 27415 96637 27493 96683
rect 27539 96637 27617 96683
rect 27663 96637 27741 96683
rect 27787 96637 27865 96683
rect 27911 96637 27989 96683
rect 28035 96637 28113 96683
rect 28159 96637 28237 96683
rect 28283 96637 28361 96683
rect 28407 96637 28485 96683
rect 28531 96637 28609 96683
rect 28655 96637 28733 96683
rect 28779 96637 28857 96683
rect 28903 96637 28981 96683
rect 29027 96637 29105 96683
rect 29151 96637 29229 96683
rect 29275 96637 29353 96683
rect 29399 96637 29477 96683
rect 29523 96637 29601 96683
rect 29647 96637 29725 96683
rect 29771 96637 29849 96683
rect 29895 96637 29973 96683
rect 30019 96637 30097 96683
rect 30143 96637 30221 96683
rect 30267 96637 30345 96683
rect 30391 96637 30469 96683
rect 30515 96637 30593 96683
rect 30639 96637 30717 96683
rect 30763 96637 30841 96683
rect 30887 96637 30965 96683
rect 31011 96637 31089 96683
rect 31135 96637 31213 96683
rect 31259 96637 31337 96683
rect 31383 96637 31461 96683
rect 31507 96637 31585 96683
rect 31631 96637 31709 96683
rect 31755 96637 31833 96683
rect 31879 96637 31957 96683
rect 32003 96637 32081 96683
rect 32127 96637 32205 96683
rect 32251 96637 32329 96683
rect 32375 96637 32453 96683
rect 32499 96637 32577 96683
rect 32623 96637 32701 96683
rect 32747 96637 32825 96683
rect 32871 96637 32949 96683
rect 32995 96637 33073 96683
rect 33119 96637 33197 96683
rect 33243 96637 33321 96683
rect 33367 96637 33445 96683
rect 33491 96637 33569 96683
rect 33615 96637 33693 96683
rect 33739 96637 33817 96683
rect 33863 96637 33941 96683
rect 33987 96637 34065 96683
rect 34111 96637 34189 96683
rect 34235 96637 34313 96683
rect 34359 96637 34437 96683
rect 34483 96637 34561 96683
rect 34607 96637 34685 96683
rect 34731 96637 34809 96683
rect 34855 96637 34933 96683
rect 34979 96637 35057 96683
rect 35103 96637 35181 96683
rect 35227 96637 35305 96683
rect 35351 96637 35429 96683
rect 35475 96637 35553 96683
rect 35599 96637 35677 96683
rect 35723 96637 35801 96683
rect 35847 96637 35925 96683
rect 35971 96637 36049 96683
rect 36095 96637 36173 96683
rect 36219 96637 36297 96683
rect 36343 96637 36421 96683
rect 36467 96637 36545 96683
rect 36591 96637 36669 96683
rect 36715 96637 36793 96683
rect 36839 96637 36917 96683
rect 36963 96637 37041 96683
rect 37087 96637 37165 96683
rect 37211 96637 37289 96683
rect 37335 96637 37413 96683
rect 37459 96637 37537 96683
rect 37583 96637 37661 96683
rect 37707 96637 37785 96683
rect 37831 96637 37909 96683
rect 37955 96637 38033 96683
rect 38079 96637 38157 96683
rect 38203 96637 38281 96683
rect 38327 96637 38405 96683
rect 38451 96637 38529 96683
rect 38575 96637 38653 96683
rect 38699 96637 38777 96683
rect 38823 96637 38901 96683
rect 38947 96637 39025 96683
rect 39071 96637 39149 96683
rect 39195 96637 39273 96683
rect 39319 96637 39397 96683
rect 39443 96637 39521 96683
rect 39567 96637 39645 96683
rect 39691 96637 39769 96683
rect 39815 96637 39893 96683
rect 39939 96637 40017 96683
rect 40063 96637 40141 96683
rect 40187 96637 40265 96683
rect 40311 96637 40389 96683
rect 40435 96637 40513 96683
rect 40559 96637 40637 96683
rect 40683 96637 40761 96683
rect 40807 96637 40885 96683
rect 40931 96637 41009 96683
rect 41055 96637 41133 96683
rect 41179 96637 41257 96683
rect 41303 96637 41381 96683
rect 41427 96637 41505 96683
rect 41551 96637 41629 96683
rect 41675 96637 41753 96683
rect 41799 96637 41877 96683
rect 41923 96637 42001 96683
rect 42047 96637 42125 96683
rect 42171 96637 42249 96683
rect 42295 96637 42373 96683
rect 42419 96637 42497 96683
rect 42543 96637 42621 96683
rect 42667 96637 42745 96683
rect 42791 96637 42869 96683
rect 42915 96637 42993 96683
rect 43039 96637 43117 96683
rect 43163 96637 43241 96683
rect 43287 96637 43365 96683
rect 43411 96637 43489 96683
rect 43535 96637 43613 96683
rect 43659 96637 43737 96683
rect 43783 96637 43861 96683
rect 43907 96637 43985 96683
rect 44031 96637 44109 96683
rect 44155 96637 44233 96683
rect 44279 96637 44357 96683
rect 44403 96637 44481 96683
rect 44527 96637 44605 96683
rect 44651 96637 44729 96683
rect 44775 96637 44853 96683
rect 44899 96637 44977 96683
rect 45023 96637 45101 96683
rect 45147 96637 45225 96683
rect 45271 96637 45349 96683
rect 45395 96637 45473 96683
rect 45519 96637 45597 96683
rect 45643 96637 45721 96683
rect 45767 96637 45845 96683
rect 45891 96637 45969 96683
rect 46015 96637 46093 96683
rect 46139 96637 46217 96683
rect 46263 96637 46341 96683
rect 46387 96637 46465 96683
rect 46511 96637 46589 96683
rect 46635 96637 46713 96683
rect 46759 96637 46837 96683
rect 46883 96637 46961 96683
rect 47007 96637 47085 96683
rect 47131 96637 47209 96683
rect 47255 96637 47333 96683
rect 47379 96637 47457 96683
rect 47503 96637 47581 96683
rect 47627 96637 47705 96683
rect 47751 96637 47829 96683
rect 47875 96637 47953 96683
rect 47999 96637 48077 96683
rect 48123 96637 48201 96683
rect 48247 96637 48325 96683
rect 48371 96637 48449 96683
rect 48495 96637 48573 96683
rect 48619 96637 48697 96683
rect 48743 96637 48821 96683
rect 48867 96637 48945 96683
rect 48991 96637 49069 96683
rect 49115 96637 49193 96683
rect 49239 96637 49317 96683
rect 49363 96637 49441 96683
rect 49487 96637 49565 96683
rect 49611 96637 49689 96683
rect 49735 96637 49813 96683
rect 49859 96637 49937 96683
rect 49983 96637 50061 96683
rect 50107 96637 50185 96683
rect 50231 96637 50309 96683
rect 50355 96637 50433 96683
rect 50479 96637 50557 96683
rect 50603 96637 50681 96683
rect 50727 96637 50805 96683
rect 50851 96637 50929 96683
rect 50975 96637 51053 96683
rect 51099 96637 51177 96683
rect 51223 96637 51301 96683
rect 51347 96637 51425 96683
rect 51471 96637 51549 96683
rect 51595 96637 51673 96683
rect 51719 96637 51797 96683
rect 51843 96637 51921 96683
rect 51967 96637 52045 96683
rect 52091 96637 52169 96683
rect 52215 96637 52293 96683
rect 52339 96637 52417 96683
rect 52463 96637 52541 96683
rect 52587 96637 52665 96683
rect 52711 96637 52789 96683
rect 52835 96637 52913 96683
rect 52959 96637 53037 96683
rect 53083 96637 53161 96683
rect 53207 96637 53285 96683
rect 53331 96637 53409 96683
rect 53455 96637 53533 96683
rect 53579 96637 53657 96683
rect 53703 96637 53781 96683
rect 53827 96637 53905 96683
rect 53951 96637 54029 96683
rect 54075 96637 54153 96683
rect 54199 96637 54277 96683
rect 54323 96637 54401 96683
rect 54447 96637 54525 96683
rect 54571 96637 54649 96683
rect 54695 96637 54773 96683
rect 54819 96637 54897 96683
rect 54943 96637 55021 96683
rect 55067 96637 55145 96683
rect 55191 96637 55269 96683
rect 55315 96637 55393 96683
rect 55439 96637 55517 96683
rect 55563 96637 55641 96683
rect 55687 96637 55765 96683
rect 55811 96637 55889 96683
rect 55935 96637 56013 96683
rect 56059 96637 56137 96683
rect 56183 96637 56261 96683
rect 56307 96637 56385 96683
rect 56431 96637 56509 96683
rect 56555 96637 56633 96683
rect 56679 96637 56757 96683
rect 56803 96637 56881 96683
rect 56927 96637 57005 96683
rect 57051 96637 57129 96683
rect 57175 96637 57253 96683
rect 57299 96637 57377 96683
rect 57423 96637 57501 96683
rect 57547 96637 57625 96683
rect 57671 96637 57749 96683
rect 57795 96637 57873 96683
rect 57919 96637 57997 96683
rect 58043 96637 58121 96683
rect 58167 96637 58245 96683
rect 58291 96637 58369 96683
rect 58415 96637 58493 96683
rect 58539 96637 58617 96683
rect 58663 96637 58741 96683
rect 58787 96637 58865 96683
rect 58911 96637 58989 96683
rect 59035 96637 59113 96683
rect 59159 96637 59237 96683
rect 59283 96637 59361 96683
rect 59407 96637 59485 96683
rect 59531 96637 59609 96683
rect 59655 96637 59733 96683
rect 59779 96637 59857 96683
rect 59903 96637 59981 96683
rect 60027 96637 60105 96683
rect 60151 96637 60229 96683
rect 60275 96637 60353 96683
rect 60399 96637 60477 96683
rect 60523 96637 60601 96683
rect 60647 96637 60725 96683
rect 60771 96637 60849 96683
rect 60895 96637 60973 96683
rect 61019 96637 61097 96683
rect 61143 96637 61221 96683
rect 61267 96637 61345 96683
rect 61391 96637 61469 96683
rect 61515 96637 61593 96683
rect 61639 96637 61717 96683
rect 61763 96637 61841 96683
rect 61887 96637 61965 96683
rect 62011 96637 62089 96683
rect 62135 96637 62213 96683
rect 62259 96637 62337 96683
rect 62383 96637 62461 96683
rect 62507 96637 62585 96683
rect 62631 96637 62709 96683
rect 62755 96637 62833 96683
rect 62879 96637 62957 96683
rect 63003 96637 63081 96683
rect 63127 96637 63205 96683
rect 63251 96637 63329 96683
rect 63375 96637 63453 96683
rect 63499 96637 63577 96683
rect 63623 96637 63701 96683
rect 63747 96637 63825 96683
rect 63871 96637 63949 96683
rect 63995 96637 64073 96683
rect 64119 96637 64197 96683
rect 64243 96637 64321 96683
rect 64367 96637 64445 96683
rect 64491 96637 64569 96683
rect 64615 96637 64693 96683
rect 64739 96637 64817 96683
rect 64863 96637 64941 96683
rect 64987 96637 65065 96683
rect 65111 96637 65189 96683
rect 65235 96637 65313 96683
rect 65359 96637 65437 96683
rect 65483 96637 65561 96683
rect 65607 96637 65685 96683
rect 65731 96637 65809 96683
rect 65855 96637 65933 96683
rect 65979 96637 66057 96683
rect 66103 96637 66181 96683
rect 66227 96637 66305 96683
rect 66351 96637 66429 96683
rect 66475 96637 66553 96683
rect 66599 96637 66677 96683
rect 66723 96637 66801 96683
rect 66847 96637 66925 96683
rect 66971 96637 67049 96683
rect 67095 96637 67173 96683
rect 67219 96637 67297 96683
rect 67343 96637 67421 96683
rect 67467 96637 67545 96683
rect 67591 96637 67669 96683
rect 67715 96637 67793 96683
rect 67839 96637 67917 96683
rect 67963 96637 68041 96683
rect 68087 96637 68165 96683
rect 68211 96637 68289 96683
rect 68335 96637 68413 96683
rect 68459 96637 68537 96683
rect 68583 96637 68661 96683
rect 68707 96637 68785 96683
rect 68831 96637 68909 96683
rect 68955 96637 69033 96683
rect 69079 96637 69157 96683
rect 69203 96637 69281 96683
rect 69327 96637 69405 96683
rect 69451 96637 69529 96683
rect 69575 96637 69653 96683
rect 69699 96637 69777 96683
rect 69823 96637 69901 96683
rect 69947 96637 70025 96683
rect 70071 96637 70149 96683
rect 70195 96637 70273 96683
rect 70319 96637 70397 96683
rect 70443 96637 70521 96683
rect 70567 96637 70645 96683
rect 70691 96637 70769 96683
rect 70815 96637 70893 96683
rect 70939 96637 71017 96683
rect 71063 96637 71141 96683
rect 71187 96637 71265 96683
rect 71311 96637 71389 96683
rect 71435 96637 71513 96683
rect 71559 96637 71637 96683
rect 71683 96637 71761 96683
rect 71807 96637 71885 96683
rect 71931 96637 72009 96683
rect 72055 96637 72133 96683
rect 72179 96637 72257 96683
rect 72303 96637 72381 96683
rect 72427 96637 72505 96683
rect 72551 96637 72629 96683
rect 72675 96637 72753 96683
rect 72799 96637 72877 96683
rect 72923 96637 73001 96683
rect 73047 96637 73125 96683
rect 73171 96637 73249 96683
rect 73295 96637 73373 96683
rect 73419 96637 73497 96683
rect 73543 96637 73621 96683
rect 73667 96637 73745 96683
rect 73791 96637 73869 96683
rect 73915 96637 73993 96683
rect 74039 96637 74117 96683
rect 74163 96637 74241 96683
rect 74287 96637 74365 96683
rect 74411 96637 74489 96683
rect 74535 96637 74613 96683
rect 74659 96637 74737 96683
rect 74783 96637 74861 96683
rect 74907 96637 74985 96683
rect 75031 96637 75109 96683
rect 75155 96637 75233 96683
rect 75279 96637 75357 96683
rect 75403 96637 75481 96683
rect 75527 96637 75605 96683
rect 75651 96637 75729 96683
rect 75775 96637 75853 96683
rect 75899 96637 75977 96683
rect 76023 96637 76101 96683
rect 76147 96637 76225 96683
rect 76271 96637 76349 96683
rect 76395 96637 76473 96683
rect 76519 96637 76597 96683
rect 76643 96637 76721 96683
rect 76767 96637 76845 96683
rect 76891 96637 76969 96683
rect 77015 96637 77093 96683
rect 77139 96637 77217 96683
rect 77263 96637 77341 96683
rect 77387 96637 77465 96683
rect 77511 96637 77589 96683
rect 77635 96637 77713 96683
rect 77759 96637 77837 96683
rect 77883 96637 77961 96683
rect 78007 96637 78085 96683
rect 78131 96637 78209 96683
rect 78255 96637 78333 96683
rect 78379 96637 78457 96683
rect 78503 96637 78581 96683
rect 78627 96637 78705 96683
rect 78751 96637 78829 96683
rect 78875 96637 78953 96683
rect 78999 96637 79077 96683
rect 79123 96637 79201 96683
rect 79247 96637 79325 96683
rect 79371 96637 79449 96683
rect 79495 96637 79573 96683
rect 79619 96637 79697 96683
rect 79743 96637 79821 96683
rect 79867 96637 79945 96683
rect 79991 96637 80069 96683
rect 80115 96637 80193 96683
rect 80239 96637 80317 96683
rect 80363 96637 80441 96683
rect 80487 96637 80565 96683
rect 80611 96637 80689 96683
rect 80735 96637 80813 96683
rect 80859 96637 80937 96683
rect 80983 96637 81061 96683
rect 81107 96637 81185 96683
rect 81231 96637 81309 96683
rect 81355 96637 81433 96683
rect 81479 96637 81557 96683
rect 81603 96637 81681 96683
rect 81727 96637 81805 96683
rect 81851 96637 81929 96683
rect 81975 96637 82053 96683
rect 82099 96637 82177 96683
rect 82223 96637 82301 96683
rect 82347 96637 82425 96683
rect 82471 96637 82549 96683
rect 82595 96637 82673 96683
rect 82719 96637 82797 96683
rect 82843 96637 82921 96683
rect 82967 96637 83045 96683
rect 83091 96637 83169 96683
rect 83215 96637 83293 96683
rect 83339 96637 83417 96683
rect 83463 96637 83541 96683
rect 83587 96637 83665 96683
rect 83711 96637 83789 96683
rect 83835 96637 83913 96683
rect 83959 96637 84037 96683
rect 84083 96637 84161 96683
rect 84207 96637 84285 96683
rect 84331 96637 84409 96683
rect 84455 96637 84533 96683
rect 84579 96637 84657 96683
rect 84703 96637 84781 96683
rect 84827 96637 84905 96683
rect 84951 96637 85029 96683
rect 85075 96637 85153 96683
rect 85199 96637 85277 96683
rect 85323 96637 85401 96683
rect 85447 96637 85525 96683
rect 85571 96637 85649 96683
rect 85695 96637 85816 96683
rect 70 96559 85816 96637
rect 70 96513 89 96559
rect 135 96513 213 96559
rect 259 96513 337 96559
rect 383 96513 461 96559
rect 507 96513 585 96559
rect 631 96513 709 96559
rect 755 96513 833 96559
rect 879 96513 957 96559
rect 1003 96513 1081 96559
rect 1127 96513 1205 96559
rect 1251 96513 1329 96559
rect 1375 96513 1453 96559
rect 1499 96513 1577 96559
rect 1623 96513 1701 96559
rect 1747 96513 1825 96559
rect 1871 96513 1949 96559
rect 1995 96513 2073 96559
rect 2119 96513 2197 96559
rect 2243 96513 2321 96559
rect 2367 96513 2445 96559
rect 2491 96513 2569 96559
rect 2615 96513 2693 96559
rect 2739 96513 2817 96559
rect 2863 96513 2941 96559
rect 2987 96513 3065 96559
rect 3111 96513 3189 96559
rect 3235 96513 3313 96559
rect 3359 96513 3437 96559
rect 3483 96513 3561 96559
rect 3607 96513 3685 96559
rect 3731 96513 3809 96559
rect 3855 96513 3933 96559
rect 3979 96513 4057 96559
rect 4103 96513 4181 96559
rect 4227 96513 4305 96559
rect 4351 96513 4429 96559
rect 4475 96513 4553 96559
rect 4599 96513 4677 96559
rect 4723 96513 4801 96559
rect 4847 96513 4925 96559
rect 4971 96513 5049 96559
rect 5095 96513 5173 96559
rect 5219 96513 5297 96559
rect 5343 96513 5421 96559
rect 5467 96513 5545 96559
rect 5591 96513 5669 96559
rect 5715 96513 5793 96559
rect 5839 96513 5917 96559
rect 5963 96513 6041 96559
rect 6087 96513 6165 96559
rect 6211 96513 6289 96559
rect 6335 96513 6413 96559
rect 6459 96513 6537 96559
rect 6583 96513 6661 96559
rect 6707 96513 6785 96559
rect 6831 96513 6909 96559
rect 6955 96513 7033 96559
rect 7079 96513 7157 96559
rect 7203 96513 7281 96559
rect 7327 96513 7405 96559
rect 7451 96513 7529 96559
rect 7575 96513 7653 96559
rect 7699 96513 7777 96559
rect 7823 96513 7901 96559
rect 7947 96513 8025 96559
rect 8071 96513 8149 96559
rect 8195 96513 8273 96559
rect 8319 96513 8397 96559
rect 8443 96513 8521 96559
rect 8567 96513 8645 96559
rect 8691 96513 8769 96559
rect 8815 96513 8893 96559
rect 8939 96513 9017 96559
rect 9063 96513 9141 96559
rect 9187 96513 9265 96559
rect 9311 96513 9389 96559
rect 9435 96513 9513 96559
rect 9559 96513 9637 96559
rect 9683 96513 9761 96559
rect 9807 96513 9885 96559
rect 9931 96513 10009 96559
rect 10055 96513 10133 96559
rect 10179 96513 10257 96559
rect 10303 96513 10381 96559
rect 10427 96513 10505 96559
rect 10551 96513 10629 96559
rect 10675 96513 10753 96559
rect 10799 96513 10877 96559
rect 10923 96513 11001 96559
rect 11047 96513 11125 96559
rect 11171 96513 11249 96559
rect 11295 96513 11373 96559
rect 11419 96513 11497 96559
rect 11543 96513 11621 96559
rect 11667 96513 11745 96559
rect 11791 96513 11869 96559
rect 11915 96513 11993 96559
rect 12039 96513 12117 96559
rect 12163 96513 12241 96559
rect 12287 96513 12365 96559
rect 12411 96513 12489 96559
rect 12535 96513 12613 96559
rect 12659 96513 12737 96559
rect 12783 96513 12861 96559
rect 12907 96513 12985 96559
rect 13031 96513 13109 96559
rect 13155 96513 13233 96559
rect 13279 96513 13357 96559
rect 13403 96513 13481 96559
rect 13527 96513 13605 96559
rect 13651 96513 13729 96559
rect 13775 96513 13853 96559
rect 13899 96513 13977 96559
rect 14023 96513 14101 96559
rect 14147 96513 14225 96559
rect 14271 96513 14349 96559
rect 14395 96513 14473 96559
rect 14519 96513 14597 96559
rect 14643 96513 14721 96559
rect 14767 96513 14845 96559
rect 14891 96513 14969 96559
rect 15015 96513 15093 96559
rect 15139 96513 15217 96559
rect 15263 96513 15341 96559
rect 15387 96513 15465 96559
rect 15511 96513 15589 96559
rect 15635 96513 15713 96559
rect 15759 96513 15837 96559
rect 15883 96513 15961 96559
rect 16007 96513 16085 96559
rect 16131 96513 16209 96559
rect 16255 96513 16333 96559
rect 16379 96513 16457 96559
rect 16503 96513 16581 96559
rect 16627 96513 16705 96559
rect 16751 96513 16829 96559
rect 16875 96513 16953 96559
rect 16999 96513 17077 96559
rect 17123 96513 17201 96559
rect 17247 96513 17325 96559
rect 17371 96513 17449 96559
rect 17495 96513 17573 96559
rect 17619 96513 17697 96559
rect 17743 96513 17821 96559
rect 17867 96513 17945 96559
rect 17991 96513 18069 96559
rect 18115 96513 18193 96559
rect 18239 96513 18317 96559
rect 18363 96513 18441 96559
rect 18487 96513 18565 96559
rect 18611 96513 18689 96559
rect 18735 96513 18813 96559
rect 18859 96513 18937 96559
rect 18983 96513 19061 96559
rect 19107 96513 19185 96559
rect 19231 96513 19309 96559
rect 19355 96513 19433 96559
rect 19479 96513 19557 96559
rect 19603 96513 19681 96559
rect 19727 96513 19805 96559
rect 19851 96513 19929 96559
rect 19975 96513 20053 96559
rect 20099 96513 20177 96559
rect 20223 96513 20301 96559
rect 20347 96513 20425 96559
rect 20471 96513 20549 96559
rect 20595 96513 20673 96559
rect 20719 96513 20797 96559
rect 20843 96513 20921 96559
rect 20967 96513 21045 96559
rect 21091 96513 21169 96559
rect 21215 96513 21293 96559
rect 21339 96513 21417 96559
rect 21463 96513 21541 96559
rect 21587 96513 21665 96559
rect 21711 96513 21789 96559
rect 21835 96513 21913 96559
rect 21959 96513 22037 96559
rect 22083 96513 22161 96559
rect 22207 96513 22285 96559
rect 22331 96513 22409 96559
rect 22455 96513 22533 96559
rect 22579 96513 22657 96559
rect 22703 96513 22781 96559
rect 22827 96513 22905 96559
rect 22951 96513 23029 96559
rect 23075 96513 23153 96559
rect 23199 96513 23277 96559
rect 23323 96513 23401 96559
rect 23447 96513 23525 96559
rect 23571 96513 23649 96559
rect 23695 96513 23773 96559
rect 23819 96513 23897 96559
rect 23943 96513 24021 96559
rect 24067 96513 24145 96559
rect 24191 96513 24269 96559
rect 24315 96513 24393 96559
rect 24439 96513 24517 96559
rect 24563 96513 24641 96559
rect 24687 96513 24765 96559
rect 24811 96513 24889 96559
rect 24935 96513 25013 96559
rect 25059 96513 25137 96559
rect 25183 96513 25261 96559
rect 25307 96513 25385 96559
rect 25431 96513 25509 96559
rect 25555 96513 25633 96559
rect 25679 96513 25757 96559
rect 25803 96513 25881 96559
rect 25927 96513 26005 96559
rect 26051 96513 26129 96559
rect 26175 96513 26253 96559
rect 26299 96513 26377 96559
rect 26423 96513 26501 96559
rect 26547 96513 26625 96559
rect 26671 96513 26749 96559
rect 26795 96513 26873 96559
rect 26919 96513 26997 96559
rect 27043 96513 27121 96559
rect 27167 96513 27245 96559
rect 27291 96513 27369 96559
rect 27415 96513 27493 96559
rect 27539 96513 27617 96559
rect 27663 96513 27741 96559
rect 27787 96513 27865 96559
rect 27911 96513 27989 96559
rect 28035 96513 28113 96559
rect 28159 96513 28237 96559
rect 28283 96513 28361 96559
rect 28407 96513 28485 96559
rect 28531 96513 28609 96559
rect 28655 96513 28733 96559
rect 28779 96513 28857 96559
rect 28903 96513 28981 96559
rect 29027 96513 29105 96559
rect 29151 96513 29229 96559
rect 29275 96513 29353 96559
rect 29399 96513 29477 96559
rect 29523 96513 29601 96559
rect 29647 96513 29725 96559
rect 29771 96513 29849 96559
rect 29895 96513 29973 96559
rect 30019 96513 30097 96559
rect 30143 96513 30221 96559
rect 30267 96513 30345 96559
rect 30391 96513 30469 96559
rect 30515 96513 30593 96559
rect 30639 96513 30717 96559
rect 30763 96513 30841 96559
rect 30887 96513 30965 96559
rect 31011 96513 31089 96559
rect 31135 96513 31213 96559
rect 31259 96513 31337 96559
rect 31383 96513 31461 96559
rect 31507 96513 31585 96559
rect 31631 96513 31709 96559
rect 31755 96513 31833 96559
rect 31879 96513 31957 96559
rect 32003 96513 32081 96559
rect 32127 96513 32205 96559
rect 32251 96513 32329 96559
rect 32375 96513 32453 96559
rect 32499 96513 32577 96559
rect 32623 96513 32701 96559
rect 32747 96513 32825 96559
rect 32871 96513 32949 96559
rect 32995 96513 33073 96559
rect 33119 96513 33197 96559
rect 33243 96513 33321 96559
rect 33367 96513 33445 96559
rect 33491 96513 33569 96559
rect 33615 96513 33693 96559
rect 33739 96513 33817 96559
rect 33863 96513 33941 96559
rect 33987 96513 34065 96559
rect 34111 96513 34189 96559
rect 34235 96513 34313 96559
rect 34359 96513 34437 96559
rect 34483 96513 34561 96559
rect 34607 96513 34685 96559
rect 34731 96513 34809 96559
rect 34855 96513 34933 96559
rect 34979 96513 35057 96559
rect 35103 96513 35181 96559
rect 35227 96513 35305 96559
rect 35351 96513 35429 96559
rect 35475 96513 35553 96559
rect 35599 96513 35677 96559
rect 35723 96513 35801 96559
rect 35847 96513 35925 96559
rect 35971 96513 36049 96559
rect 36095 96513 36173 96559
rect 36219 96513 36297 96559
rect 36343 96513 36421 96559
rect 36467 96513 36545 96559
rect 36591 96513 36669 96559
rect 36715 96513 36793 96559
rect 36839 96513 36917 96559
rect 36963 96513 37041 96559
rect 37087 96513 37165 96559
rect 37211 96513 37289 96559
rect 37335 96513 37413 96559
rect 37459 96513 37537 96559
rect 37583 96513 37661 96559
rect 37707 96513 37785 96559
rect 37831 96513 37909 96559
rect 37955 96513 38033 96559
rect 38079 96513 38157 96559
rect 38203 96513 38281 96559
rect 38327 96513 38405 96559
rect 38451 96513 38529 96559
rect 38575 96513 38653 96559
rect 38699 96513 38777 96559
rect 38823 96513 38901 96559
rect 38947 96513 39025 96559
rect 39071 96513 39149 96559
rect 39195 96513 39273 96559
rect 39319 96513 39397 96559
rect 39443 96513 39521 96559
rect 39567 96513 39645 96559
rect 39691 96513 39769 96559
rect 39815 96513 39893 96559
rect 39939 96513 40017 96559
rect 40063 96513 40141 96559
rect 40187 96513 40265 96559
rect 40311 96513 40389 96559
rect 40435 96513 40513 96559
rect 40559 96513 40637 96559
rect 40683 96513 40761 96559
rect 40807 96513 40885 96559
rect 40931 96513 41009 96559
rect 41055 96513 41133 96559
rect 41179 96513 41257 96559
rect 41303 96513 41381 96559
rect 41427 96513 41505 96559
rect 41551 96513 41629 96559
rect 41675 96513 41753 96559
rect 41799 96513 41877 96559
rect 41923 96513 42001 96559
rect 42047 96513 42125 96559
rect 42171 96513 42249 96559
rect 42295 96513 42373 96559
rect 42419 96513 42497 96559
rect 42543 96513 42621 96559
rect 42667 96513 42745 96559
rect 42791 96513 42869 96559
rect 42915 96513 42993 96559
rect 43039 96513 43117 96559
rect 43163 96513 43241 96559
rect 43287 96513 43365 96559
rect 43411 96513 43489 96559
rect 43535 96513 43613 96559
rect 43659 96513 43737 96559
rect 43783 96513 43861 96559
rect 43907 96513 43985 96559
rect 44031 96513 44109 96559
rect 44155 96513 44233 96559
rect 44279 96513 44357 96559
rect 44403 96513 44481 96559
rect 44527 96513 44605 96559
rect 44651 96513 44729 96559
rect 44775 96513 44853 96559
rect 44899 96513 44977 96559
rect 45023 96513 45101 96559
rect 45147 96513 45225 96559
rect 45271 96513 45349 96559
rect 45395 96513 45473 96559
rect 45519 96513 45597 96559
rect 45643 96513 45721 96559
rect 45767 96513 45845 96559
rect 45891 96513 45969 96559
rect 46015 96513 46093 96559
rect 46139 96513 46217 96559
rect 46263 96513 46341 96559
rect 46387 96513 46465 96559
rect 46511 96513 46589 96559
rect 46635 96513 46713 96559
rect 46759 96513 46837 96559
rect 46883 96513 46961 96559
rect 47007 96513 47085 96559
rect 47131 96513 47209 96559
rect 47255 96513 47333 96559
rect 47379 96513 47457 96559
rect 47503 96513 47581 96559
rect 47627 96513 47705 96559
rect 47751 96513 47829 96559
rect 47875 96513 47953 96559
rect 47999 96513 48077 96559
rect 48123 96513 48201 96559
rect 48247 96513 48325 96559
rect 48371 96513 48449 96559
rect 48495 96513 48573 96559
rect 48619 96513 48697 96559
rect 48743 96513 48821 96559
rect 48867 96513 48945 96559
rect 48991 96513 49069 96559
rect 49115 96513 49193 96559
rect 49239 96513 49317 96559
rect 49363 96513 49441 96559
rect 49487 96513 49565 96559
rect 49611 96513 49689 96559
rect 49735 96513 49813 96559
rect 49859 96513 49937 96559
rect 49983 96513 50061 96559
rect 50107 96513 50185 96559
rect 50231 96513 50309 96559
rect 50355 96513 50433 96559
rect 50479 96513 50557 96559
rect 50603 96513 50681 96559
rect 50727 96513 50805 96559
rect 50851 96513 50929 96559
rect 50975 96513 51053 96559
rect 51099 96513 51177 96559
rect 51223 96513 51301 96559
rect 51347 96513 51425 96559
rect 51471 96513 51549 96559
rect 51595 96513 51673 96559
rect 51719 96513 51797 96559
rect 51843 96513 51921 96559
rect 51967 96513 52045 96559
rect 52091 96513 52169 96559
rect 52215 96513 52293 96559
rect 52339 96513 52417 96559
rect 52463 96513 52541 96559
rect 52587 96513 52665 96559
rect 52711 96513 52789 96559
rect 52835 96513 52913 96559
rect 52959 96513 53037 96559
rect 53083 96513 53161 96559
rect 53207 96513 53285 96559
rect 53331 96513 53409 96559
rect 53455 96513 53533 96559
rect 53579 96513 53657 96559
rect 53703 96513 53781 96559
rect 53827 96513 53905 96559
rect 53951 96513 54029 96559
rect 54075 96513 54153 96559
rect 54199 96513 54277 96559
rect 54323 96513 54401 96559
rect 54447 96513 54525 96559
rect 54571 96513 54649 96559
rect 54695 96513 54773 96559
rect 54819 96513 54897 96559
rect 54943 96513 55021 96559
rect 55067 96513 55145 96559
rect 55191 96513 55269 96559
rect 55315 96513 55393 96559
rect 55439 96513 55517 96559
rect 55563 96513 55641 96559
rect 55687 96513 55765 96559
rect 55811 96513 55889 96559
rect 55935 96513 56013 96559
rect 56059 96513 56137 96559
rect 56183 96513 56261 96559
rect 56307 96513 56385 96559
rect 56431 96513 56509 96559
rect 56555 96513 56633 96559
rect 56679 96513 56757 96559
rect 56803 96513 56881 96559
rect 56927 96513 57005 96559
rect 57051 96513 57129 96559
rect 57175 96513 57253 96559
rect 57299 96513 57377 96559
rect 57423 96513 57501 96559
rect 57547 96513 57625 96559
rect 57671 96513 57749 96559
rect 57795 96513 57873 96559
rect 57919 96513 57997 96559
rect 58043 96513 58121 96559
rect 58167 96513 58245 96559
rect 58291 96513 58369 96559
rect 58415 96513 58493 96559
rect 58539 96513 58617 96559
rect 58663 96513 58741 96559
rect 58787 96513 58865 96559
rect 58911 96513 58989 96559
rect 59035 96513 59113 96559
rect 59159 96513 59237 96559
rect 59283 96513 59361 96559
rect 59407 96513 59485 96559
rect 59531 96513 59609 96559
rect 59655 96513 59733 96559
rect 59779 96513 59857 96559
rect 59903 96513 59981 96559
rect 60027 96513 60105 96559
rect 60151 96513 60229 96559
rect 60275 96513 60353 96559
rect 60399 96513 60477 96559
rect 60523 96513 60601 96559
rect 60647 96513 60725 96559
rect 60771 96513 60849 96559
rect 60895 96513 60973 96559
rect 61019 96513 61097 96559
rect 61143 96513 61221 96559
rect 61267 96513 61345 96559
rect 61391 96513 61469 96559
rect 61515 96513 61593 96559
rect 61639 96513 61717 96559
rect 61763 96513 61841 96559
rect 61887 96513 61965 96559
rect 62011 96513 62089 96559
rect 62135 96513 62213 96559
rect 62259 96513 62337 96559
rect 62383 96513 62461 96559
rect 62507 96513 62585 96559
rect 62631 96513 62709 96559
rect 62755 96513 62833 96559
rect 62879 96513 62957 96559
rect 63003 96513 63081 96559
rect 63127 96513 63205 96559
rect 63251 96513 63329 96559
rect 63375 96513 63453 96559
rect 63499 96513 63577 96559
rect 63623 96513 63701 96559
rect 63747 96513 63825 96559
rect 63871 96513 63949 96559
rect 63995 96513 64073 96559
rect 64119 96513 64197 96559
rect 64243 96513 64321 96559
rect 64367 96513 64445 96559
rect 64491 96513 64569 96559
rect 64615 96513 64693 96559
rect 64739 96513 64817 96559
rect 64863 96513 64941 96559
rect 64987 96513 65065 96559
rect 65111 96513 65189 96559
rect 65235 96513 65313 96559
rect 65359 96513 65437 96559
rect 65483 96513 65561 96559
rect 65607 96513 65685 96559
rect 65731 96513 65809 96559
rect 65855 96513 65933 96559
rect 65979 96513 66057 96559
rect 66103 96513 66181 96559
rect 66227 96513 66305 96559
rect 66351 96513 66429 96559
rect 66475 96513 66553 96559
rect 66599 96513 66677 96559
rect 66723 96513 66801 96559
rect 66847 96513 66925 96559
rect 66971 96513 67049 96559
rect 67095 96513 67173 96559
rect 67219 96513 67297 96559
rect 67343 96513 67421 96559
rect 67467 96513 67545 96559
rect 67591 96513 67669 96559
rect 67715 96513 67793 96559
rect 67839 96513 67917 96559
rect 67963 96513 68041 96559
rect 68087 96513 68165 96559
rect 68211 96513 68289 96559
rect 68335 96513 68413 96559
rect 68459 96513 68537 96559
rect 68583 96513 68661 96559
rect 68707 96513 68785 96559
rect 68831 96513 68909 96559
rect 68955 96513 69033 96559
rect 69079 96513 69157 96559
rect 69203 96513 69281 96559
rect 69327 96513 69405 96559
rect 69451 96513 69529 96559
rect 69575 96513 69653 96559
rect 69699 96513 69777 96559
rect 69823 96513 69901 96559
rect 69947 96513 70025 96559
rect 70071 96513 70149 96559
rect 70195 96513 70273 96559
rect 70319 96513 70397 96559
rect 70443 96513 70521 96559
rect 70567 96513 70645 96559
rect 70691 96513 70769 96559
rect 70815 96513 70893 96559
rect 70939 96513 71017 96559
rect 71063 96513 71141 96559
rect 71187 96513 71265 96559
rect 71311 96513 71389 96559
rect 71435 96513 71513 96559
rect 71559 96513 71637 96559
rect 71683 96513 71761 96559
rect 71807 96513 71885 96559
rect 71931 96513 72009 96559
rect 72055 96513 72133 96559
rect 72179 96513 72257 96559
rect 72303 96513 72381 96559
rect 72427 96513 72505 96559
rect 72551 96513 72629 96559
rect 72675 96513 72753 96559
rect 72799 96513 72877 96559
rect 72923 96513 73001 96559
rect 73047 96513 73125 96559
rect 73171 96513 73249 96559
rect 73295 96513 73373 96559
rect 73419 96513 73497 96559
rect 73543 96513 73621 96559
rect 73667 96513 73745 96559
rect 73791 96513 73869 96559
rect 73915 96513 73993 96559
rect 74039 96513 74117 96559
rect 74163 96513 74241 96559
rect 74287 96513 74365 96559
rect 74411 96513 74489 96559
rect 74535 96513 74613 96559
rect 74659 96513 74737 96559
rect 74783 96513 74861 96559
rect 74907 96513 74985 96559
rect 75031 96513 75109 96559
rect 75155 96513 75233 96559
rect 75279 96513 75357 96559
rect 75403 96513 75481 96559
rect 75527 96513 75605 96559
rect 75651 96513 75729 96559
rect 75775 96513 75853 96559
rect 75899 96513 75977 96559
rect 76023 96513 76101 96559
rect 76147 96513 76225 96559
rect 76271 96513 76349 96559
rect 76395 96513 76473 96559
rect 76519 96513 76597 96559
rect 76643 96513 76721 96559
rect 76767 96513 76845 96559
rect 76891 96513 76969 96559
rect 77015 96513 77093 96559
rect 77139 96513 77217 96559
rect 77263 96513 77341 96559
rect 77387 96513 77465 96559
rect 77511 96513 77589 96559
rect 77635 96513 77713 96559
rect 77759 96513 77837 96559
rect 77883 96513 77961 96559
rect 78007 96513 78085 96559
rect 78131 96513 78209 96559
rect 78255 96513 78333 96559
rect 78379 96513 78457 96559
rect 78503 96513 78581 96559
rect 78627 96513 78705 96559
rect 78751 96513 78829 96559
rect 78875 96513 78953 96559
rect 78999 96513 79077 96559
rect 79123 96513 79201 96559
rect 79247 96513 79325 96559
rect 79371 96513 79449 96559
rect 79495 96513 79573 96559
rect 79619 96513 79697 96559
rect 79743 96513 79821 96559
rect 79867 96513 79945 96559
rect 79991 96513 80069 96559
rect 80115 96513 80193 96559
rect 80239 96513 80317 96559
rect 80363 96513 80441 96559
rect 80487 96513 80565 96559
rect 80611 96513 80689 96559
rect 80735 96513 80813 96559
rect 80859 96513 80937 96559
rect 80983 96513 81061 96559
rect 81107 96513 81185 96559
rect 81231 96513 81309 96559
rect 81355 96513 81433 96559
rect 81479 96513 81557 96559
rect 81603 96513 81681 96559
rect 81727 96513 81805 96559
rect 81851 96513 81929 96559
rect 81975 96513 82053 96559
rect 82099 96513 82177 96559
rect 82223 96513 82301 96559
rect 82347 96513 82425 96559
rect 82471 96513 82549 96559
rect 82595 96513 82673 96559
rect 82719 96513 82797 96559
rect 82843 96513 82921 96559
rect 82967 96513 83045 96559
rect 83091 96513 83169 96559
rect 83215 96513 83293 96559
rect 83339 96513 83417 96559
rect 83463 96513 83541 96559
rect 83587 96513 83665 96559
rect 83711 96513 83789 96559
rect 83835 96513 83913 96559
rect 83959 96513 84037 96559
rect 84083 96513 84161 96559
rect 84207 96513 84285 96559
rect 84331 96513 84409 96559
rect 84455 96513 84533 96559
rect 84579 96513 84657 96559
rect 84703 96513 84781 96559
rect 84827 96513 84905 96559
rect 84951 96513 85029 96559
rect 85075 96513 85153 96559
rect 85199 96513 85277 96559
rect 85323 96513 85401 96559
rect 85447 96513 85525 96559
rect 85571 96513 85649 96559
rect 85695 96513 85816 96559
rect 70 96435 85816 96513
rect 70 96389 89 96435
rect 135 96389 213 96435
rect 259 96389 337 96435
rect 383 96389 461 96435
rect 507 96389 585 96435
rect 631 96389 709 96435
rect 755 96389 833 96435
rect 879 96389 957 96435
rect 1003 96389 1081 96435
rect 1127 96389 1205 96435
rect 1251 96389 1329 96435
rect 1375 96389 1453 96435
rect 1499 96389 1577 96435
rect 1623 96389 1701 96435
rect 1747 96389 1825 96435
rect 1871 96389 1949 96435
rect 1995 96389 2073 96435
rect 2119 96389 2197 96435
rect 2243 96389 2321 96435
rect 2367 96389 2445 96435
rect 2491 96389 2569 96435
rect 2615 96389 2693 96435
rect 2739 96389 2817 96435
rect 2863 96389 2941 96435
rect 2987 96389 3065 96435
rect 3111 96389 3189 96435
rect 3235 96389 3313 96435
rect 3359 96389 3437 96435
rect 3483 96389 3561 96435
rect 3607 96389 3685 96435
rect 3731 96389 3809 96435
rect 3855 96389 3933 96435
rect 3979 96389 4057 96435
rect 4103 96389 4181 96435
rect 4227 96389 4305 96435
rect 4351 96389 4429 96435
rect 4475 96389 4553 96435
rect 4599 96389 4677 96435
rect 4723 96389 4801 96435
rect 4847 96389 4925 96435
rect 4971 96389 5049 96435
rect 5095 96389 5173 96435
rect 5219 96389 5297 96435
rect 5343 96389 5421 96435
rect 5467 96389 5545 96435
rect 5591 96389 5669 96435
rect 5715 96389 5793 96435
rect 5839 96389 5917 96435
rect 5963 96389 6041 96435
rect 6087 96389 6165 96435
rect 6211 96389 6289 96435
rect 6335 96389 6413 96435
rect 6459 96389 6537 96435
rect 6583 96389 6661 96435
rect 6707 96389 6785 96435
rect 6831 96389 6909 96435
rect 6955 96389 7033 96435
rect 7079 96389 7157 96435
rect 7203 96389 7281 96435
rect 7327 96389 7405 96435
rect 7451 96389 7529 96435
rect 7575 96389 7653 96435
rect 7699 96389 7777 96435
rect 7823 96389 7901 96435
rect 7947 96389 8025 96435
rect 8071 96389 8149 96435
rect 8195 96389 8273 96435
rect 8319 96389 8397 96435
rect 8443 96389 8521 96435
rect 8567 96389 8645 96435
rect 8691 96389 8769 96435
rect 8815 96389 8893 96435
rect 8939 96389 9017 96435
rect 9063 96389 9141 96435
rect 9187 96389 9265 96435
rect 9311 96389 9389 96435
rect 9435 96389 9513 96435
rect 9559 96389 9637 96435
rect 9683 96389 9761 96435
rect 9807 96389 9885 96435
rect 9931 96389 10009 96435
rect 10055 96389 10133 96435
rect 10179 96389 10257 96435
rect 10303 96389 10381 96435
rect 10427 96389 10505 96435
rect 10551 96389 10629 96435
rect 10675 96389 10753 96435
rect 10799 96389 10877 96435
rect 10923 96389 11001 96435
rect 11047 96389 11125 96435
rect 11171 96389 11249 96435
rect 11295 96389 11373 96435
rect 11419 96389 11497 96435
rect 11543 96389 11621 96435
rect 11667 96389 11745 96435
rect 11791 96389 11869 96435
rect 11915 96389 11993 96435
rect 12039 96389 12117 96435
rect 12163 96389 12241 96435
rect 12287 96389 12365 96435
rect 12411 96389 12489 96435
rect 12535 96389 12613 96435
rect 12659 96389 12737 96435
rect 12783 96389 12861 96435
rect 12907 96389 12985 96435
rect 13031 96389 13109 96435
rect 13155 96389 13233 96435
rect 13279 96389 13357 96435
rect 13403 96389 13481 96435
rect 13527 96389 13605 96435
rect 13651 96389 13729 96435
rect 13775 96389 13853 96435
rect 13899 96389 13977 96435
rect 14023 96389 14101 96435
rect 14147 96389 14225 96435
rect 14271 96389 14349 96435
rect 14395 96389 14473 96435
rect 14519 96389 14597 96435
rect 14643 96389 14721 96435
rect 14767 96389 14845 96435
rect 14891 96389 14969 96435
rect 15015 96389 15093 96435
rect 15139 96389 15217 96435
rect 15263 96389 15341 96435
rect 15387 96389 15465 96435
rect 15511 96389 15589 96435
rect 15635 96389 15713 96435
rect 15759 96389 15837 96435
rect 15883 96389 15961 96435
rect 16007 96389 16085 96435
rect 16131 96389 16209 96435
rect 16255 96389 16333 96435
rect 16379 96389 16457 96435
rect 16503 96389 16581 96435
rect 16627 96389 16705 96435
rect 16751 96389 16829 96435
rect 16875 96389 16953 96435
rect 16999 96389 17077 96435
rect 17123 96389 17201 96435
rect 17247 96389 17325 96435
rect 17371 96389 17449 96435
rect 17495 96389 17573 96435
rect 17619 96389 17697 96435
rect 17743 96389 17821 96435
rect 17867 96389 17945 96435
rect 17991 96389 18069 96435
rect 18115 96389 18193 96435
rect 18239 96389 18317 96435
rect 18363 96389 18441 96435
rect 18487 96389 18565 96435
rect 18611 96389 18689 96435
rect 18735 96389 18813 96435
rect 18859 96389 18937 96435
rect 18983 96389 19061 96435
rect 19107 96389 19185 96435
rect 19231 96389 19309 96435
rect 19355 96389 19433 96435
rect 19479 96389 19557 96435
rect 19603 96389 19681 96435
rect 19727 96389 19805 96435
rect 19851 96389 19929 96435
rect 19975 96389 20053 96435
rect 20099 96389 20177 96435
rect 20223 96389 20301 96435
rect 20347 96389 20425 96435
rect 20471 96389 20549 96435
rect 20595 96389 20673 96435
rect 20719 96389 20797 96435
rect 20843 96389 20921 96435
rect 20967 96389 21045 96435
rect 21091 96389 21169 96435
rect 21215 96389 21293 96435
rect 21339 96389 21417 96435
rect 21463 96389 21541 96435
rect 21587 96389 21665 96435
rect 21711 96389 21789 96435
rect 21835 96389 21913 96435
rect 21959 96389 22037 96435
rect 22083 96389 22161 96435
rect 22207 96389 22285 96435
rect 22331 96389 22409 96435
rect 22455 96389 22533 96435
rect 22579 96389 22657 96435
rect 22703 96389 22781 96435
rect 22827 96389 22905 96435
rect 22951 96389 23029 96435
rect 23075 96389 23153 96435
rect 23199 96389 23277 96435
rect 23323 96389 23401 96435
rect 23447 96389 23525 96435
rect 23571 96389 23649 96435
rect 23695 96389 23773 96435
rect 23819 96389 23897 96435
rect 23943 96389 24021 96435
rect 24067 96389 24145 96435
rect 24191 96389 24269 96435
rect 24315 96389 24393 96435
rect 24439 96389 24517 96435
rect 24563 96389 24641 96435
rect 24687 96389 24765 96435
rect 24811 96389 24889 96435
rect 24935 96389 25013 96435
rect 25059 96389 25137 96435
rect 25183 96389 25261 96435
rect 25307 96389 25385 96435
rect 25431 96389 25509 96435
rect 25555 96389 25633 96435
rect 25679 96389 25757 96435
rect 25803 96389 25881 96435
rect 25927 96389 26005 96435
rect 26051 96389 26129 96435
rect 26175 96389 26253 96435
rect 26299 96389 26377 96435
rect 26423 96389 26501 96435
rect 26547 96389 26625 96435
rect 26671 96389 26749 96435
rect 26795 96389 26873 96435
rect 26919 96389 26997 96435
rect 27043 96389 27121 96435
rect 27167 96389 27245 96435
rect 27291 96389 27369 96435
rect 27415 96389 27493 96435
rect 27539 96389 27617 96435
rect 27663 96389 27741 96435
rect 27787 96389 27865 96435
rect 27911 96389 27989 96435
rect 28035 96389 28113 96435
rect 28159 96389 28237 96435
rect 28283 96389 28361 96435
rect 28407 96389 28485 96435
rect 28531 96389 28609 96435
rect 28655 96389 28733 96435
rect 28779 96389 28857 96435
rect 28903 96389 28981 96435
rect 29027 96389 29105 96435
rect 29151 96389 29229 96435
rect 29275 96389 29353 96435
rect 29399 96389 29477 96435
rect 29523 96389 29601 96435
rect 29647 96389 29725 96435
rect 29771 96389 29849 96435
rect 29895 96389 29973 96435
rect 30019 96389 30097 96435
rect 30143 96389 30221 96435
rect 30267 96389 30345 96435
rect 30391 96389 30469 96435
rect 30515 96389 30593 96435
rect 30639 96389 30717 96435
rect 30763 96389 30841 96435
rect 30887 96389 30965 96435
rect 31011 96389 31089 96435
rect 31135 96389 31213 96435
rect 31259 96389 31337 96435
rect 31383 96389 31461 96435
rect 31507 96389 31585 96435
rect 31631 96389 31709 96435
rect 31755 96389 31833 96435
rect 31879 96389 31957 96435
rect 32003 96389 32081 96435
rect 32127 96389 32205 96435
rect 32251 96389 32329 96435
rect 32375 96389 32453 96435
rect 32499 96389 32577 96435
rect 32623 96389 32701 96435
rect 32747 96389 32825 96435
rect 32871 96389 32949 96435
rect 32995 96389 33073 96435
rect 33119 96389 33197 96435
rect 33243 96389 33321 96435
rect 33367 96389 33445 96435
rect 33491 96389 33569 96435
rect 33615 96389 33693 96435
rect 33739 96389 33817 96435
rect 33863 96389 33941 96435
rect 33987 96389 34065 96435
rect 34111 96389 34189 96435
rect 34235 96389 34313 96435
rect 34359 96389 34437 96435
rect 34483 96389 34561 96435
rect 34607 96389 34685 96435
rect 34731 96389 34809 96435
rect 34855 96389 34933 96435
rect 34979 96389 35057 96435
rect 35103 96389 35181 96435
rect 35227 96389 35305 96435
rect 35351 96389 35429 96435
rect 35475 96389 35553 96435
rect 35599 96389 35677 96435
rect 35723 96389 35801 96435
rect 35847 96389 35925 96435
rect 35971 96389 36049 96435
rect 36095 96389 36173 96435
rect 36219 96389 36297 96435
rect 36343 96389 36421 96435
rect 36467 96389 36545 96435
rect 36591 96389 36669 96435
rect 36715 96389 36793 96435
rect 36839 96389 36917 96435
rect 36963 96389 37041 96435
rect 37087 96389 37165 96435
rect 37211 96389 37289 96435
rect 37335 96389 37413 96435
rect 37459 96389 37537 96435
rect 37583 96389 37661 96435
rect 37707 96389 37785 96435
rect 37831 96389 37909 96435
rect 37955 96389 38033 96435
rect 38079 96389 38157 96435
rect 38203 96389 38281 96435
rect 38327 96389 38405 96435
rect 38451 96389 38529 96435
rect 38575 96389 38653 96435
rect 38699 96389 38777 96435
rect 38823 96389 38901 96435
rect 38947 96389 39025 96435
rect 39071 96389 39149 96435
rect 39195 96389 39273 96435
rect 39319 96389 39397 96435
rect 39443 96389 39521 96435
rect 39567 96389 39645 96435
rect 39691 96389 39769 96435
rect 39815 96389 39893 96435
rect 39939 96389 40017 96435
rect 40063 96389 40141 96435
rect 40187 96389 40265 96435
rect 40311 96389 40389 96435
rect 40435 96389 40513 96435
rect 40559 96389 40637 96435
rect 40683 96389 40761 96435
rect 40807 96389 40885 96435
rect 40931 96389 41009 96435
rect 41055 96389 41133 96435
rect 41179 96389 41257 96435
rect 41303 96389 41381 96435
rect 41427 96389 41505 96435
rect 41551 96389 41629 96435
rect 41675 96389 41753 96435
rect 41799 96389 41877 96435
rect 41923 96389 42001 96435
rect 42047 96389 42125 96435
rect 42171 96389 42249 96435
rect 42295 96389 42373 96435
rect 42419 96389 42497 96435
rect 42543 96389 42621 96435
rect 42667 96389 42745 96435
rect 42791 96389 42869 96435
rect 42915 96389 42993 96435
rect 43039 96389 43117 96435
rect 43163 96389 43241 96435
rect 43287 96389 43365 96435
rect 43411 96389 43489 96435
rect 43535 96389 43613 96435
rect 43659 96389 43737 96435
rect 43783 96389 43861 96435
rect 43907 96389 43985 96435
rect 44031 96389 44109 96435
rect 44155 96389 44233 96435
rect 44279 96389 44357 96435
rect 44403 96389 44481 96435
rect 44527 96389 44605 96435
rect 44651 96389 44729 96435
rect 44775 96389 44853 96435
rect 44899 96389 44977 96435
rect 45023 96389 45101 96435
rect 45147 96389 45225 96435
rect 45271 96389 45349 96435
rect 45395 96389 45473 96435
rect 45519 96389 45597 96435
rect 45643 96389 45721 96435
rect 45767 96389 45845 96435
rect 45891 96389 45969 96435
rect 46015 96389 46093 96435
rect 46139 96389 46217 96435
rect 46263 96389 46341 96435
rect 46387 96389 46465 96435
rect 46511 96389 46589 96435
rect 46635 96389 46713 96435
rect 46759 96389 46837 96435
rect 46883 96389 46961 96435
rect 47007 96389 47085 96435
rect 47131 96389 47209 96435
rect 47255 96389 47333 96435
rect 47379 96389 47457 96435
rect 47503 96389 47581 96435
rect 47627 96389 47705 96435
rect 47751 96389 47829 96435
rect 47875 96389 47953 96435
rect 47999 96389 48077 96435
rect 48123 96389 48201 96435
rect 48247 96389 48325 96435
rect 48371 96389 48449 96435
rect 48495 96389 48573 96435
rect 48619 96389 48697 96435
rect 48743 96389 48821 96435
rect 48867 96389 48945 96435
rect 48991 96389 49069 96435
rect 49115 96389 49193 96435
rect 49239 96389 49317 96435
rect 49363 96389 49441 96435
rect 49487 96389 49565 96435
rect 49611 96389 49689 96435
rect 49735 96389 49813 96435
rect 49859 96389 49937 96435
rect 49983 96389 50061 96435
rect 50107 96389 50185 96435
rect 50231 96389 50309 96435
rect 50355 96389 50433 96435
rect 50479 96389 50557 96435
rect 50603 96389 50681 96435
rect 50727 96389 50805 96435
rect 50851 96389 50929 96435
rect 50975 96389 51053 96435
rect 51099 96389 51177 96435
rect 51223 96389 51301 96435
rect 51347 96389 51425 96435
rect 51471 96389 51549 96435
rect 51595 96389 51673 96435
rect 51719 96389 51797 96435
rect 51843 96389 51921 96435
rect 51967 96389 52045 96435
rect 52091 96389 52169 96435
rect 52215 96389 52293 96435
rect 52339 96389 52417 96435
rect 52463 96389 52541 96435
rect 52587 96389 52665 96435
rect 52711 96389 52789 96435
rect 52835 96389 52913 96435
rect 52959 96389 53037 96435
rect 53083 96389 53161 96435
rect 53207 96389 53285 96435
rect 53331 96389 53409 96435
rect 53455 96389 53533 96435
rect 53579 96389 53657 96435
rect 53703 96389 53781 96435
rect 53827 96389 53905 96435
rect 53951 96389 54029 96435
rect 54075 96389 54153 96435
rect 54199 96389 54277 96435
rect 54323 96389 54401 96435
rect 54447 96389 54525 96435
rect 54571 96389 54649 96435
rect 54695 96389 54773 96435
rect 54819 96389 54897 96435
rect 54943 96389 55021 96435
rect 55067 96389 55145 96435
rect 55191 96389 55269 96435
rect 55315 96389 55393 96435
rect 55439 96389 55517 96435
rect 55563 96389 55641 96435
rect 55687 96389 55765 96435
rect 55811 96389 55889 96435
rect 55935 96389 56013 96435
rect 56059 96389 56137 96435
rect 56183 96389 56261 96435
rect 56307 96389 56385 96435
rect 56431 96389 56509 96435
rect 56555 96389 56633 96435
rect 56679 96389 56757 96435
rect 56803 96389 56881 96435
rect 56927 96389 57005 96435
rect 57051 96389 57129 96435
rect 57175 96389 57253 96435
rect 57299 96389 57377 96435
rect 57423 96389 57501 96435
rect 57547 96389 57625 96435
rect 57671 96389 57749 96435
rect 57795 96389 57873 96435
rect 57919 96389 57997 96435
rect 58043 96389 58121 96435
rect 58167 96389 58245 96435
rect 58291 96389 58369 96435
rect 58415 96389 58493 96435
rect 58539 96389 58617 96435
rect 58663 96389 58741 96435
rect 58787 96389 58865 96435
rect 58911 96389 58989 96435
rect 59035 96389 59113 96435
rect 59159 96389 59237 96435
rect 59283 96389 59361 96435
rect 59407 96389 59485 96435
rect 59531 96389 59609 96435
rect 59655 96389 59733 96435
rect 59779 96389 59857 96435
rect 59903 96389 59981 96435
rect 60027 96389 60105 96435
rect 60151 96389 60229 96435
rect 60275 96389 60353 96435
rect 60399 96389 60477 96435
rect 60523 96389 60601 96435
rect 60647 96389 60725 96435
rect 60771 96389 60849 96435
rect 60895 96389 60973 96435
rect 61019 96389 61097 96435
rect 61143 96389 61221 96435
rect 61267 96389 61345 96435
rect 61391 96389 61469 96435
rect 61515 96389 61593 96435
rect 61639 96389 61717 96435
rect 61763 96389 61841 96435
rect 61887 96389 61965 96435
rect 62011 96389 62089 96435
rect 62135 96389 62213 96435
rect 62259 96389 62337 96435
rect 62383 96389 62461 96435
rect 62507 96389 62585 96435
rect 62631 96389 62709 96435
rect 62755 96389 62833 96435
rect 62879 96389 62957 96435
rect 63003 96389 63081 96435
rect 63127 96389 63205 96435
rect 63251 96389 63329 96435
rect 63375 96389 63453 96435
rect 63499 96389 63577 96435
rect 63623 96389 63701 96435
rect 63747 96389 63825 96435
rect 63871 96389 63949 96435
rect 63995 96389 64073 96435
rect 64119 96389 64197 96435
rect 64243 96389 64321 96435
rect 64367 96389 64445 96435
rect 64491 96389 64569 96435
rect 64615 96389 64693 96435
rect 64739 96389 64817 96435
rect 64863 96389 64941 96435
rect 64987 96389 65065 96435
rect 65111 96389 65189 96435
rect 65235 96389 65313 96435
rect 65359 96389 65437 96435
rect 65483 96389 65561 96435
rect 65607 96389 65685 96435
rect 65731 96389 65809 96435
rect 65855 96389 65933 96435
rect 65979 96389 66057 96435
rect 66103 96389 66181 96435
rect 66227 96389 66305 96435
rect 66351 96389 66429 96435
rect 66475 96389 66553 96435
rect 66599 96389 66677 96435
rect 66723 96389 66801 96435
rect 66847 96389 66925 96435
rect 66971 96389 67049 96435
rect 67095 96389 67173 96435
rect 67219 96389 67297 96435
rect 67343 96389 67421 96435
rect 67467 96389 67545 96435
rect 67591 96389 67669 96435
rect 67715 96389 67793 96435
rect 67839 96389 67917 96435
rect 67963 96389 68041 96435
rect 68087 96389 68165 96435
rect 68211 96389 68289 96435
rect 68335 96389 68413 96435
rect 68459 96389 68537 96435
rect 68583 96389 68661 96435
rect 68707 96389 68785 96435
rect 68831 96389 68909 96435
rect 68955 96389 69033 96435
rect 69079 96389 69157 96435
rect 69203 96389 69281 96435
rect 69327 96389 69405 96435
rect 69451 96389 69529 96435
rect 69575 96389 69653 96435
rect 69699 96389 69777 96435
rect 69823 96389 69901 96435
rect 69947 96389 70025 96435
rect 70071 96389 70149 96435
rect 70195 96389 70273 96435
rect 70319 96389 70397 96435
rect 70443 96389 70521 96435
rect 70567 96389 70645 96435
rect 70691 96389 70769 96435
rect 70815 96389 70893 96435
rect 70939 96389 71017 96435
rect 71063 96389 71141 96435
rect 71187 96389 71265 96435
rect 71311 96389 71389 96435
rect 71435 96389 71513 96435
rect 71559 96389 71637 96435
rect 71683 96389 71761 96435
rect 71807 96389 71885 96435
rect 71931 96389 72009 96435
rect 72055 96389 72133 96435
rect 72179 96389 72257 96435
rect 72303 96389 72381 96435
rect 72427 96389 72505 96435
rect 72551 96389 72629 96435
rect 72675 96389 72753 96435
rect 72799 96389 72877 96435
rect 72923 96389 73001 96435
rect 73047 96389 73125 96435
rect 73171 96389 73249 96435
rect 73295 96389 73373 96435
rect 73419 96389 73497 96435
rect 73543 96389 73621 96435
rect 73667 96389 73745 96435
rect 73791 96389 73869 96435
rect 73915 96389 73993 96435
rect 74039 96389 74117 96435
rect 74163 96389 74241 96435
rect 74287 96389 74365 96435
rect 74411 96389 74489 96435
rect 74535 96389 74613 96435
rect 74659 96389 74737 96435
rect 74783 96389 74861 96435
rect 74907 96389 74985 96435
rect 75031 96389 75109 96435
rect 75155 96389 75233 96435
rect 75279 96389 75357 96435
rect 75403 96389 75481 96435
rect 75527 96389 75605 96435
rect 75651 96389 75729 96435
rect 75775 96389 75853 96435
rect 75899 96389 75977 96435
rect 76023 96389 76101 96435
rect 76147 96389 76225 96435
rect 76271 96389 76349 96435
rect 76395 96389 76473 96435
rect 76519 96389 76597 96435
rect 76643 96389 76721 96435
rect 76767 96389 76845 96435
rect 76891 96389 76969 96435
rect 77015 96389 77093 96435
rect 77139 96389 77217 96435
rect 77263 96389 77341 96435
rect 77387 96389 77465 96435
rect 77511 96389 77589 96435
rect 77635 96389 77713 96435
rect 77759 96389 77837 96435
rect 77883 96389 77961 96435
rect 78007 96389 78085 96435
rect 78131 96389 78209 96435
rect 78255 96389 78333 96435
rect 78379 96389 78457 96435
rect 78503 96389 78581 96435
rect 78627 96389 78705 96435
rect 78751 96389 78829 96435
rect 78875 96389 78953 96435
rect 78999 96389 79077 96435
rect 79123 96389 79201 96435
rect 79247 96389 79325 96435
rect 79371 96389 79449 96435
rect 79495 96389 79573 96435
rect 79619 96389 79697 96435
rect 79743 96389 79821 96435
rect 79867 96389 79945 96435
rect 79991 96389 80069 96435
rect 80115 96389 80193 96435
rect 80239 96389 80317 96435
rect 80363 96389 80441 96435
rect 80487 96389 80565 96435
rect 80611 96389 80689 96435
rect 80735 96389 80813 96435
rect 80859 96389 80937 96435
rect 80983 96389 81061 96435
rect 81107 96389 81185 96435
rect 81231 96389 81309 96435
rect 81355 96389 81433 96435
rect 81479 96389 81557 96435
rect 81603 96389 81681 96435
rect 81727 96389 81805 96435
rect 81851 96389 81929 96435
rect 81975 96389 82053 96435
rect 82099 96389 82177 96435
rect 82223 96389 82301 96435
rect 82347 96389 82425 96435
rect 82471 96389 82549 96435
rect 82595 96389 82673 96435
rect 82719 96389 82797 96435
rect 82843 96389 82921 96435
rect 82967 96389 83045 96435
rect 83091 96389 83169 96435
rect 83215 96389 83293 96435
rect 83339 96389 83417 96435
rect 83463 96389 83541 96435
rect 83587 96389 83665 96435
rect 83711 96389 83789 96435
rect 83835 96389 83913 96435
rect 83959 96389 84037 96435
rect 84083 96389 84161 96435
rect 84207 96389 84285 96435
rect 84331 96389 84409 96435
rect 84455 96389 84533 96435
rect 84579 96389 84657 96435
rect 84703 96389 84781 96435
rect 84827 96389 84905 96435
rect 84951 96389 85029 96435
rect 85075 96389 85153 96435
rect 85199 96389 85277 96435
rect 85323 96389 85401 96435
rect 85447 96389 85525 96435
rect 85571 96389 85649 96435
rect 85695 96389 85816 96435
rect 70 96311 85816 96389
rect 70 96265 89 96311
rect 135 96265 213 96311
rect 259 96265 337 96311
rect 383 96265 461 96311
rect 507 96265 585 96311
rect 631 96265 709 96311
rect 755 96265 833 96311
rect 879 96265 957 96311
rect 1003 96265 1081 96311
rect 1127 96265 1205 96311
rect 1251 96265 1329 96311
rect 1375 96265 1453 96311
rect 1499 96265 1577 96311
rect 1623 96265 1701 96311
rect 1747 96265 1825 96311
rect 1871 96265 1949 96311
rect 1995 96265 2073 96311
rect 2119 96265 2197 96311
rect 2243 96265 2321 96311
rect 2367 96265 2445 96311
rect 2491 96265 2569 96311
rect 2615 96265 2693 96311
rect 2739 96265 2817 96311
rect 2863 96265 2941 96311
rect 2987 96265 3065 96311
rect 3111 96265 3189 96311
rect 3235 96265 3313 96311
rect 3359 96265 3437 96311
rect 3483 96265 3561 96311
rect 3607 96265 3685 96311
rect 3731 96265 3809 96311
rect 3855 96265 3933 96311
rect 3979 96265 4057 96311
rect 4103 96265 4181 96311
rect 4227 96265 4305 96311
rect 4351 96265 4429 96311
rect 4475 96265 4553 96311
rect 4599 96265 4677 96311
rect 4723 96265 4801 96311
rect 4847 96265 4925 96311
rect 4971 96265 5049 96311
rect 5095 96265 5173 96311
rect 5219 96265 5297 96311
rect 5343 96265 5421 96311
rect 5467 96265 5545 96311
rect 5591 96265 5669 96311
rect 5715 96265 5793 96311
rect 5839 96265 5917 96311
rect 5963 96265 6041 96311
rect 6087 96265 6165 96311
rect 6211 96265 6289 96311
rect 6335 96265 6413 96311
rect 6459 96265 6537 96311
rect 6583 96265 6661 96311
rect 6707 96265 6785 96311
rect 6831 96265 6909 96311
rect 6955 96265 7033 96311
rect 7079 96265 7157 96311
rect 7203 96265 7281 96311
rect 7327 96265 7405 96311
rect 7451 96265 7529 96311
rect 7575 96265 7653 96311
rect 7699 96265 7777 96311
rect 7823 96265 7901 96311
rect 7947 96265 8025 96311
rect 8071 96265 8149 96311
rect 8195 96265 8273 96311
rect 8319 96265 8397 96311
rect 8443 96265 8521 96311
rect 8567 96265 8645 96311
rect 8691 96265 8769 96311
rect 8815 96265 8893 96311
rect 8939 96265 9017 96311
rect 9063 96265 9141 96311
rect 9187 96265 9265 96311
rect 9311 96265 9389 96311
rect 9435 96265 9513 96311
rect 9559 96265 9637 96311
rect 9683 96265 9761 96311
rect 9807 96265 9885 96311
rect 9931 96265 10009 96311
rect 10055 96265 10133 96311
rect 10179 96265 10257 96311
rect 10303 96265 10381 96311
rect 10427 96265 10505 96311
rect 10551 96265 10629 96311
rect 10675 96265 10753 96311
rect 10799 96265 10877 96311
rect 10923 96265 11001 96311
rect 11047 96265 11125 96311
rect 11171 96265 11249 96311
rect 11295 96265 11373 96311
rect 11419 96265 11497 96311
rect 11543 96265 11621 96311
rect 11667 96265 11745 96311
rect 11791 96265 11869 96311
rect 11915 96265 11993 96311
rect 12039 96265 12117 96311
rect 12163 96265 12241 96311
rect 12287 96265 12365 96311
rect 12411 96265 12489 96311
rect 12535 96265 12613 96311
rect 12659 96265 12737 96311
rect 12783 96265 12861 96311
rect 12907 96265 12985 96311
rect 13031 96265 13109 96311
rect 13155 96265 13233 96311
rect 13279 96265 13357 96311
rect 13403 96265 13481 96311
rect 13527 96265 13605 96311
rect 13651 96265 13729 96311
rect 13775 96265 13853 96311
rect 13899 96265 13977 96311
rect 14023 96265 14101 96311
rect 14147 96265 14225 96311
rect 14271 96265 14349 96311
rect 14395 96265 14473 96311
rect 14519 96265 14597 96311
rect 14643 96265 14721 96311
rect 14767 96265 14845 96311
rect 14891 96265 14969 96311
rect 15015 96265 15093 96311
rect 15139 96265 15217 96311
rect 15263 96265 15341 96311
rect 15387 96265 15465 96311
rect 15511 96265 15589 96311
rect 15635 96265 15713 96311
rect 15759 96265 15837 96311
rect 15883 96265 15961 96311
rect 16007 96265 16085 96311
rect 16131 96265 16209 96311
rect 16255 96265 16333 96311
rect 16379 96265 16457 96311
rect 16503 96265 16581 96311
rect 16627 96265 16705 96311
rect 16751 96265 16829 96311
rect 16875 96265 16953 96311
rect 16999 96265 17077 96311
rect 17123 96265 17201 96311
rect 17247 96265 17325 96311
rect 17371 96265 17449 96311
rect 17495 96265 17573 96311
rect 17619 96265 17697 96311
rect 17743 96265 17821 96311
rect 17867 96265 17945 96311
rect 17991 96265 18069 96311
rect 18115 96265 18193 96311
rect 18239 96265 18317 96311
rect 18363 96265 18441 96311
rect 18487 96265 18565 96311
rect 18611 96265 18689 96311
rect 18735 96265 18813 96311
rect 18859 96265 18937 96311
rect 18983 96265 19061 96311
rect 19107 96265 19185 96311
rect 19231 96265 19309 96311
rect 19355 96265 19433 96311
rect 19479 96265 19557 96311
rect 19603 96265 19681 96311
rect 19727 96265 19805 96311
rect 19851 96265 19929 96311
rect 19975 96265 20053 96311
rect 20099 96265 20177 96311
rect 20223 96265 20301 96311
rect 20347 96265 20425 96311
rect 20471 96265 20549 96311
rect 20595 96265 20673 96311
rect 20719 96265 20797 96311
rect 20843 96265 20921 96311
rect 20967 96265 21045 96311
rect 21091 96265 21169 96311
rect 21215 96265 21293 96311
rect 21339 96265 21417 96311
rect 21463 96265 21541 96311
rect 21587 96265 21665 96311
rect 21711 96265 21789 96311
rect 21835 96265 21913 96311
rect 21959 96265 22037 96311
rect 22083 96265 22161 96311
rect 22207 96265 22285 96311
rect 22331 96265 22409 96311
rect 22455 96265 22533 96311
rect 22579 96265 22657 96311
rect 22703 96265 22781 96311
rect 22827 96265 22905 96311
rect 22951 96265 23029 96311
rect 23075 96265 23153 96311
rect 23199 96265 23277 96311
rect 23323 96265 23401 96311
rect 23447 96265 23525 96311
rect 23571 96265 23649 96311
rect 23695 96265 23773 96311
rect 23819 96265 23897 96311
rect 23943 96265 24021 96311
rect 24067 96265 24145 96311
rect 24191 96265 24269 96311
rect 24315 96265 24393 96311
rect 24439 96265 24517 96311
rect 24563 96265 24641 96311
rect 24687 96265 24765 96311
rect 24811 96265 24889 96311
rect 24935 96265 25013 96311
rect 25059 96265 25137 96311
rect 25183 96265 25261 96311
rect 25307 96265 25385 96311
rect 25431 96265 25509 96311
rect 25555 96265 25633 96311
rect 25679 96265 25757 96311
rect 25803 96265 25881 96311
rect 25927 96265 26005 96311
rect 26051 96265 26129 96311
rect 26175 96265 26253 96311
rect 26299 96265 26377 96311
rect 26423 96265 26501 96311
rect 26547 96265 26625 96311
rect 26671 96265 26749 96311
rect 26795 96265 26873 96311
rect 26919 96265 26997 96311
rect 27043 96265 27121 96311
rect 27167 96265 27245 96311
rect 27291 96265 27369 96311
rect 27415 96265 27493 96311
rect 27539 96265 27617 96311
rect 27663 96265 27741 96311
rect 27787 96265 27865 96311
rect 27911 96265 27989 96311
rect 28035 96265 28113 96311
rect 28159 96265 28237 96311
rect 28283 96265 28361 96311
rect 28407 96265 28485 96311
rect 28531 96265 28609 96311
rect 28655 96265 28733 96311
rect 28779 96265 28857 96311
rect 28903 96265 28981 96311
rect 29027 96265 29105 96311
rect 29151 96265 29229 96311
rect 29275 96265 29353 96311
rect 29399 96265 29477 96311
rect 29523 96265 29601 96311
rect 29647 96265 29725 96311
rect 29771 96265 29849 96311
rect 29895 96265 29973 96311
rect 30019 96265 30097 96311
rect 30143 96265 30221 96311
rect 30267 96265 30345 96311
rect 30391 96265 30469 96311
rect 30515 96265 30593 96311
rect 30639 96265 30717 96311
rect 30763 96265 30841 96311
rect 30887 96265 30965 96311
rect 31011 96265 31089 96311
rect 31135 96265 31213 96311
rect 31259 96265 31337 96311
rect 31383 96265 31461 96311
rect 31507 96265 31585 96311
rect 31631 96265 31709 96311
rect 31755 96265 31833 96311
rect 31879 96265 31957 96311
rect 32003 96265 32081 96311
rect 32127 96265 32205 96311
rect 32251 96265 32329 96311
rect 32375 96265 32453 96311
rect 32499 96265 32577 96311
rect 32623 96265 32701 96311
rect 32747 96265 32825 96311
rect 32871 96265 32949 96311
rect 32995 96265 33073 96311
rect 33119 96265 33197 96311
rect 33243 96265 33321 96311
rect 33367 96265 33445 96311
rect 33491 96265 33569 96311
rect 33615 96265 33693 96311
rect 33739 96265 33817 96311
rect 33863 96265 33941 96311
rect 33987 96265 34065 96311
rect 34111 96265 34189 96311
rect 34235 96265 34313 96311
rect 34359 96265 34437 96311
rect 34483 96265 34561 96311
rect 34607 96265 34685 96311
rect 34731 96265 34809 96311
rect 34855 96265 34933 96311
rect 34979 96265 35057 96311
rect 35103 96265 35181 96311
rect 35227 96265 35305 96311
rect 35351 96265 35429 96311
rect 35475 96265 35553 96311
rect 35599 96265 35677 96311
rect 35723 96265 35801 96311
rect 35847 96265 35925 96311
rect 35971 96265 36049 96311
rect 36095 96265 36173 96311
rect 36219 96265 36297 96311
rect 36343 96265 36421 96311
rect 36467 96265 36545 96311
rect 36591 96265 36669 96311
rect 36715 96265 36793 96311
rect 36839 96265 36917 96311
rect 36963 96265 37041 96311
rect 37087 96265 37165 96311
rect 37211 96265 37289 96311
rect 37335 96265 37413 96311
rect 37459 96265 37537 96311
rect 37583 96265 37661 96311
rect 37707 96265 37785 96311
rect 37831 96265 37909 96311
rect 37955 96265 38033 96311
rect 38079 96265 38157 96311
rect 38203 96265 38281 96311
rect 38327 96265 38405 96311
rect 38451 96265 38529 96311
rect 38575 96265 38653 96311
rect 38699 96265 38777 96311
rect 38823 96265 38901 96311
rect 38947 96265 39025 96311
rect 39071 96265 39149 96311
rect 39195 96265 39273 96311
rect 39319 96265 39397 96311
rect 39443 96265 39521 96311
rect 39567 96265 39645 96311
rect 39691 96265 39769 96311
rect 39815 96265 39893 96311
rect 39939 96265 40017 96311
rect 40063 96265 40141 96311
rect 40187 96265 40265 96311
rect 40311 96265 40389 96311
rect 40435 96265 40513 96311
rect 40559 96265 40637 96311
rect 40683 96265 40761 96311
rect 40807 96265 40885 96311
rect 40931 96265 41009 96311
rect 41055 96265 41133 96311
rect 41179 96265 41257 96311
rect 41303 96265 41381 96311
rect 41427 96265 41505 96311
rect 41551 96265 41629 96311
rect 41675 96265 41753 96311
rect 41799 96265 41877 96311
rect 41923 96265 42001 96311
rect 42047 96265 42125 96311
rect 42171 96265 42249 96311
rect 42295 96265 42373 96311
rect 42419 96265 42497 96311
rect 42543 96265 42621 96311
rect 42667 96265 42745 96311
rect 42791 96265 42869 96311
rect 42915 96265 42993 96311
rect 43039 96265 43117 96311
rect 43163 96265 43241 96311
rect 43287 96265 43365 96311
rect 43411 96265 43489 96311
rect 43535 96265 43613 96311
rect 43659 96265 43737 96311
rect 43783 96265 43861 96311
rect 43907 96265 43985 96311
rect 44031 96265 44109 96311
rect 44155 96265 44233 96311
rect 44279 96265 44357 96311
rect 44403 96265 44481 96311
rect 44527 96265 44605 96311
rect 44651 96265 44729 96311
rect 44775 96265 44853 96311
rect 44899 96265 44977 96311
rect 45023 96265 45101 96311
rect 45147 96265 45225 96311
rect 45271 96265 45349 96311
rect 45395 96265 45473 96311
rect 45519 96265 45597 96311
rect 45643 96265 45721 96311
rect 45767 96265 45845 96311
rect 45891 96265 45969 96311
rect 46015 96265 46093 96311
rect 46139 96265 46217 96311
rect 46263 96265 46341 96311
rect 46387 96265 46465 96311
rect 46511 96265 46589 96311
rect 46635 96265 46713 96311
rect 46759 96265 46837 96311
rect 46883 96265 46961 96311
rect 47007 96265 47085 96311
rect 47131 96265 47209 96311
rect 47255 96265 47333 96311
rect 47379 96265 47457 96311
rect 47503 96265 47581 96311
rect 47627 96265 47705 96311
rect 47751 96265 47829 96311
rect 47875 96265 47953 96311
rect 47999 96265 48077 96311
rect 48123 96265 48201 96311
rect 48247 96265 48325 96311
rect 48371 96265 48449 96311
rect 48495 96265 48573 96311
rect 48619 96265 48697 96311
rect 48743 96265 48821 96311
rect 48867 96265 48945 96311
rect 48991 96265 49069 96311
rect 49115 96265 49193 96311
rect 49239 96265 49317 96311
rect 49363 96265 49441 96311
rect 49487 96265 49565 96311
rect 49611 96265 49689 96311
rect 49735 96265 49813 96311
rect 49859 96265 49937 96311
rect 49983 96265 50061 96311
rect 50107 96265 50185 96311
rect 50231 96265 50309 96311
rect 50355 96265 50433 96311
rect 50479 96265 50557 96311
rect 50603 96265 50681 96311
rect 50727 96265 50805 96311
rect 50851 96265 50929 96311
rect 50975 96265 51053 96311
rect 51099 96265 51177 96311
rect 51223 96265 51301 96311
rect 51347 96265 51425 96311
rect 51471 96265 51549 96311
rect 51595 96265 51673 96311
rect 51719 96265 51797 96311
rect 51843 96265 51921 96311
rect 51967 96265 52045 96311
rect 52091 96265 52169 96311
rect 52215 96265 52293 96311
rect 52339 96265 52417 96311
rect 52463 96265 52541 96311
rect 52587 96265 52665 96311
rect 52711 96265 52789 96311
rect 52835 96265 52913 96311
rect 52959 96265 53037 96311
rect 53083 96265 53161 96311
rect 53207 96265 53285 96311
rect 53331 96265 53409 96311
rect 53455 96265 53533 96311
rect 53579 96265 53657 96311
rect 53703 96265 53781 96311
rect 53827 96265 53905 96311
rect 53951 96265 54029 96311
rect 54075 96265 54153 96311
rect 54199 96265 54277 96311
rect 54323 96265 54401 96311
rect 54447 96265 54525 96311
rect 54571 96265 54649 96311
rect 54695 96265 54773 96311
rect 54819 96265 54897 96311
rect 54943 96265 55021 96311
rect 55067 96265 55145 96311
rect 55191 96265 55269 96311
rect 55315 96265 55393 96311
rect 55439 96265 55517 96311
rect 55563 96265 55641 96311
rect 55687 96265 55765 96311
rect 55811 96265 55889 96311
rect 55935 96265 56013 96311
rect 56059 96265 56137 96311
rect 56183 96265 56261 96311
rect 56307 96265 56385 96311
rect 56431 96265 56509 96311
rect 56555 96265 56633 96311
rect 56679 96265 56757 96311
rect 56803 96265 56881 96311
rect 56927 96265 57005 96311
rect 57051 96265 57129 96311
rect 57175 96265 57253 96311
rect 57299 96265 57377 96311
rect 57423 96265 57501 96311
rect 57547 96265 57625 96311
rect 57671 96265 57749 96311
rect 57795 96265 57873 96311
rect 57919 96265 57997 96311
rect 58043 96265 58121 96311
rect 58167 96265 58245 96311
rect 58291 96265 58369 96311
rect 58415 96265 58493 96311
rect 58539 96265 58617 96311
rect 58663 96265 58741 96311
rect 58787 96265 58865 96311
rect 58911 96265 58989 96311
rect 59035 96265 59113 96311
rect 59159 96265 59237 96311
rect 59283 96265 59361 96311
rect 59407 96265 59485 96311
rect 59531 96265 59609 96311
rect 59655 96265 59733 96311
rect 59779 96265 59857 96311
rect 59903 96265 59981 96311
rect 60027 96265 60105 96311
rect 60151 96265 60229 96311
rect 60275 96265 60353 96311
rect 60399 96265 60477 96311
rect 60523 96265 60601 96311
rect 60647 96265 60725 96311
rect 60771 96265 60849 96311
rect 60895 96265 60973 96311
rect 61019 96265 61097 96311
rect 61143 96265 61221 96311
rect 61267 96265 61345 96311
rect 61391 96265 61469 96311
rect 61515 96265 61593 96311
rect 61639 96265 61717 96311
rect 61763 96265 61841 96311
rect 61887 96265 61965 96311
rect 62011 96265 62089 96311
rect 62135 96265 62213 96311
rect 62259 96265 62337 96311
rect 62383 96265 62461 96311
rect 62507 96265 62585 96311
rect 62631 96265 62709 96311
rect 62755 96265 62833 96311
rect 62879 96265 62957 96311
rect 63003 96265 63081 96311
rect 63127 96265 63205 96311
rect 63251 96265 63329 96311
rect 63375 96265 63453 96311
rect 63499 96265 63577 96311
rect 63623 96265 63701 96311
rect 63747 96265 63825 96311
rect 63871 96265 63949 96311
rect 63995 96265 64073 96311
rect 64119 96265 64197 96311
rect 64243 96265 64321 96311
rect 64367 96265 64445 96311
rect 64491 96265 64569 96311
rect 64615 96265 64693 96311
rect 64739 96265 64817 96311
rect 64863 96265 64941 96311
rect 64987 96265 65065 96311
rect 65111 96265 65189 96311
rect 65235 96265 65313 96311
rect 65359 96265 65437 96311
rect 65483 96265 65561 96311
rect 65607 96265 65685 96311
rect 65731 96265 65809 96311
rect 65855 96265 65933 96311
rect 65979 96265 66057 96311
rect 66103 96265 66181 96311
rect 66227 96265 66305 96311
rect 66351 96265 66429 96311
rect 66475 96265 66553 96311
rect 66599 96265 66677 96311
rect 66723 96265 66801 96311
rect 66847 96265 66925 96311
rect 66971 96265 67049 96311
rect 67095 96265 67173 96311
rect 67219 96265 67297 96311
rect 67343 96265 67421 96311
rect 67467 96265 67545 96311
rect 67591 96265 67669 96311
rect 67715 96265 67793 96311
rect 67839 96265 67917 96311
rect 67963 96265 68041 96311
rect 68087 96265 68165 96311
rect 68211 96265 68289 96311
rect 68335 96265 68413 96311
rect 68459 96265 68537 96311
rect 68583 96265 68661 96311
rect 68707 96265 68785 96311
rect 68831 96265 68909 96311
rect 68955 96265 69033 96311
rect 69079 96265 69157 96311
rect 69203 96265 69281 96311
rect 69327 96265 69405 96311
rect 69451 96265 69529 96311
rect 69575 96265 69653 96311
rect 69699 96265 69777 96311
rect 69823 96265 69901 96311
rect 69947 96265 70025 96311
rect 70071 96265 70149 96311
rect 70195 96265 70273 96311
rect 70319 96265 70397 96311
rect 70443 96265 70521 96311
rect 70567 96265 70645 96311
rect 70691 96265 70769 96311
rect 70815 96265 70893 96311
rect 70939 96265 71017 96311
rect 71063 96265 71141 96311
rect 71187 96265 71265 96311
rect 71311 96265 71389 96311
rect 71435 96265 71513 96311
rect 71559 96265 71637 96311
rect 71683 96265 71761 96311
rect 71807 96265 71885 96311
rect 71931 96265 72009 96311
rect 72055 96265 72133 96311
rect 72179 96265 72257 96311
rect 72303 96265 72381 96311
rect 72427 96265 72505 96311
rect 72551 96265 72629 96311
rect 72675 96265 72753 96311
rect 72799 96265 72877 96311
rect 72923 96265 73001 96311
rect 73047 96265 73125 96311
rect 73171 96265 73249 96311
rect 73295 96265 73373 96311
rect 73419 96265 73497 96311
rect 73543 96265 73621 96311
rect 73667 96265 73745 96311
rect 73791 96265 73869 96311
rect 73915 96265 73993 96311
rect 74039 96265 74117 96311
rect 74163 96265 74241 96311
rect 74287 96265 74365 96311
rect 74411 96265 74489 96311
rect 74535 96265 74613 96311
rect 74659 96265 74737 96311
rect 74783 96265 74861 96311
rect 74907 96265 74985 96311
rect 75031 96265 75109 96311
rect 75155 96265 75233 96311
rect 75279 96265 75357 96311
rect 75403 96265 75481 96311
rect 75527 96265 75605 96311
rect 75651 96265 75729 96311
rect 75775 96265 75853 96311
rect 75899 96265 75977 96311
rect 76023 96265 76101 96311
rect 76147 96265 76225 96311
rect 76271 96265 76349 96311
rect 76395 96265 76473 96311
rect 76519 96265 76597 96311
rect 76643 96265 76721 96311
rect 76767 96265 76845 96311
rect 76891 96265 76969 96311
rect 77015 96265 77093 96311
rect 77139 96265 77217 96311
rect 77263 96265 77341 96311
rect 77387 96265 77465 96311
rect 77511 96265 77589 96311
rect 77635 96265 77713 96311
rect 77759 96265 77837 96311
rect 77883 96265 77961 96311
rect 78007 96265 78085 96311
rect 78131 96265 78209 96311
rect 78255 96265 78333 96311
rect 78379 96265 78457 96311
rect 78503 96265 78581 96311
rect 78627 96265 78705 96311
rect 78751 96265 78829 96311
rect 78875 96265 78953 96311
rect 78999 96265 79077 96311
rect 79123 96265 79201 96311
rect 79247 96265 79325 96311
rect 79371 96265 79449 96311
rect 79495 96265 79573 96311
rect 79619 96265 79697 96311
rect 79743 96265 79821 96311
rect 79867 96265 79945 96311
rect 79991 96265 80069 96311
rect 80115 96265 80193 96311
rect 80239 96265 80317 96311
rect 80363 96265 80441 96311
rect 80487 96265 80565 96311
rect 80611 96265 80689 96311
rect 80735 96265 80813 96311
rect 80859 96265 80937 96311
rect 80983 96265 81061 96311
rect 81107 96265 81185 96311
rect 81231 96265 81309 96311
rect 81355 96265 81433 96311
rect 81479 96265 81557 96311
rect 81603 96265 81681 96311
rect 81727 96265 81805 96311
rect 81851 96265 81929 96311
rect 81975 96265 82053 96311
rect 82099 96265 82177 96311
rect 82223 96265 82301 96311
rect 82347 96265 82425 96311
rect 82471 96265 82549 96311
rect 82595 96265 82673 96311
rect 82719 96265 82797 96311
rect 82843 96265 82921 96311
rect 82967 96265 83045 96311
rect 83091 96265 83169 96311
rect 83215 96265 83293 96311
rect 83339 96265 83417 96311
rect 83463 96265 83541 96311
rect 83587 96265 83665 96311
rect 83711 96265 83789 96311
rect 83835 96265 83913 96311
rect 83959 96265 84037 96311
rect 84083 96265 84161 96311
rect 84207 96265 84285 96311
rect 84331 96265 84409 96311
rect 84455 96265 84533 96311
rect 84579 96265 84657 96311
rect 84703 96265 84781 96311
rect 84827 96265 84905 96311
rect 84951 96265 85029 96311
rect 85075 96265 85153 96311
rect 85199 96265 85277 96311
rect 85323 96265 85401 96311
rect 85447 96265 85525 96311
rect 85571 96265 85649 96311
rect 85695 96265 85816 96311
rect 70 96246 85816 96265
rect 70 96163 454 96246
rect 70 1117 89 96163
rect 435 1117 454 96163
rect 70 1034 454 1117
rect 27097 96163 28629 96246
rect 27097 1117 27116 96163
rect 27462 96142 28629 96163
rect 27462 35996 27540 96142
rect 28386 35996 28629 96142
rect 27462 35977 28629 35996
rect 55930 96163 57389 96246
rect 55930 96142 57024 96163
rect 55930 35996 56100 96142
rect 56946 35996 57024 96142
rect 55930 35977 57024 35996
rect 27462 1117 27481 35977
rect 27521 34620 56905 34639
rect 27521 34174 27540 34620
rect 56886 34174 56905 34620
rect 27521 34155 56905 34174
rect 27097 1034 27481 1117
rect 57005 1117 57024 35977
rect 57370 1117 57389 96163
rect 57005 1034 57389 1117
rect 85432 96163 85816 96246
rect 85432 1117 85451 96163
rect 85797 1117 85816 96163
rect 85432 1034 85816 1117
rect 70 1015 85816 1034
rect 70 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85816 1015
rect 70 891 85816 969
rect 70 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85816 891
rect 70 767 85816 845
rect 70 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85816 767
rect 70 643 85816 721
rect 70 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85816 643
rect 70 578 85816 597
<< psubdiffcont >>
rect 89 96637 135 96683
rect 213 96637 259 96683
rect 337 96637 383 96683
rect 461 96637 507 96683
rect 585 96637 631 96683
rect 709 96637 755 96683
rect 833 96637 879 96683
rect 957 96637 1003 96683
rect 1081 96637 1127 96683
rect 1205 96637 1251 96683
rect 1329 96637 1375 96683
rect 1453 96637 1499 96683
rect 1577 96637 1623 96683
rect 1701 96637 1747 96683
rect 1825 96637 1871 96683
rect 1949 96637 1995 96683
rect 2073 96637 2119 96683
rect 2197 96637 2243 96683
rect 2321 96637 2367 96683
rect 2445 96637 2491 96683
rect 2569 96637 2615 96683
rect 2693 96637 2739 96683
rect 2817 96637 2863 96683
rect 2941 96637 2987 96683
rect 3065 96637 3111 96683
rect 3189 96637 3235 96683
rect 3313 96637 3359 96683
rect 3437 96637 3483 96683
rect 3561 96637 3607 96683
rect 3685 96637 3731 96683
rect 3809 96637 3855 96683
rect 3933 96637 3979 96683
rect 4057 96637 4103 96683
rect 4181 96637 4227 96683
rect 4305 96637 4351 96683
rect 4429 96637 4475 96683
rect 4553 96637 4599 96683
rect 4677 96637 4723 96683
rect 4801 96637 4847 96683
rect 4925 96637 4971 96683
rect 5049 96637 5095 96683
rect 5173 96637 5219 96683
rect 5297 96637 5343 96683
rect 5421 96637 5467 96683
rect 5545 96637 5591 96683
rect 5669 96637 5715 96683
rect 5793 96637 5839 96683
rect 5917 96637 5963 96683
rect 6041 96637 6087 96683
rect 6165 96637 6211 96683
rect 6289 96637 6335 96683
rect 6413 96637 6459 96683
rect 6537 96637 6583 96683
rect 6661 96637 6707 96683
rect 6785 96637 6831 96683
rect 6909 96637 6955 96683
rect 7033 96637 7079 96683
rect 7157 96637 7203 96683
rect 7281 96637 7327 96683
rect 7405 96637 7451 96683
rect 7529 96637 7575 96683
rect 7653 96637 7699 96683
rect 7777 96637 7823 96683
rect 7901 96637 7947 96683
rect 8025 96637 8071 96683
rect 8149 96637 8195 96683
rect 8273 96637 8319 96683
rect 8397 96637 8443 96683
rect 8521 96637 8567 96683
rect 8645 96637 8691 96683
rect 8769 96637 8815 96683
rect 8893 96637 8939 96683
rect 9017 96637 9063 96683
rect 9141 96637 9187 96683
rect 9265 96637 9311 96683
rect 9389 96637 9435 96683
rect 9513 96637 9559 96683
rect 9637 96637 9683 96683
rect 9761 96637 9807 96683
rect 9885 96637 9931 96683
rect 10009 96637 10055 96683
rect 10133 96637 10179 96683
rect 10257 96637 10303 96683
rect 10381 96637 10427 96683
rect 10505 96637 10551 96683
rect 10629 96637 10675 96683
rect 10753 96637 10799 96683
rect 10877 96637 10923 96683
rect 11001 96637 11047 96683
rect 11125 96637 11171 96683
rect 11249 96637 11295 96683
rect 11373 96637 11419 96683
rect 11497 96637 11543 96683
rect 11621 96637 11667 96683
rect 11745 96637 11791 96683
rect 11869 96637 11915 96683
rect 11993 96637 12039 96683
rect 12117 96637 12163 96683
rect 12241 96637 12287 96683
rect 12365 96637 12411 96683
rect 12489 96637 12535 96683
rect 12613 96637 12659 96683
rect 12737 96637 12783 96683
rect 12861 96637 12907 96683
rect 12985 96637 13031 96683
rect 13109 96637 13155 96683
rect 13233 96637 13279 96683
rect 13357 96637 13403 96683
rect 13481 96637 13527 96683
rect 13605 96637 13651 96683
rect 13729 96637 13775 96683
rect 13853 96637 13899 96683
rect 13977 96637 14023 96683
rect 14101 96637 14147 96683
rect 14225 96637 14271 96683
rect 14349 96637 14395 96683
rect 14473 96637 14519 96683
rect 14597 96637 14643 96683
rect 14721 96637 14767 96683
rect 14845 96637 14891 96683
rect 14969 96637 15015 96683
rect 15093 96637 15139 96683
rect 15217 96637 15263 96683
rect 15341 96637 15387 96683
rect 15465 96637 15511 96683
rect 15589 96637 15635 96683
rect 15713 96637 15759 96683
rect 15837 96637 15883 96683
rect 15961 96637 16007 96683
rect 16085 96637 16131 96683
rect 16209 96637 16255 96683
rect 16333 96637 16379 96683
rect 16457 96637 16503 96683
rect 16581 96637 16627 96683
rect 16705 96637 16751 96683
rect 16829 96637 16875 96683
rect 16953 96637 16999 96683
rect 17077 96637 17123 96683
rect 17201 96637 17247 96683
rect 17325 96637 17371 96683
rect 17449 96637 17495 96683
rect 17573 96637 17619 96683
rect 17697 96637 17743 96683
rect 17821 96637 17867 96683
rect 17945 96637 17991 96683
rect 18069 96637 18115 96683
rect 18193 96637 18239 96683
rect 18317 96637 18363 96683
rect 18441 96637 18487 96683
rect 18565 96637 18611 96683
rect 18689 96637 18735 96683
rect 18813 96637 18859 96683
rect 18937 96637 18983 96683
rect 19061 96637 19107 96683
rect 19185 96637 19231 96683
rect 19309 96637 19355 96683
rect 19433 96637 19479 96683
rect 19557 96637 19603 96683
rect 19681 96637 19727 96683
rect 19805 96637 19851 96683
rect 19929 96637 19975 96683
rect 20053 96637 20099 96683
rect 20177 96637 20223 96683
rect 20301 96637 20347 96683
rect 20425 96637 20471 96683
rect 20549 96637 20595 96683
rect 20673 96637 20719 96683
rect 20797 96637 20843 96683
rect 20921 96637 20967 96683
rect 21045 96637 21091 96683
rect 21169 96637 21215 96683
rect 21293 96637 21339 96683
rect 21417 96637 21463 96683
rect 21541 96637 21587 96683
rect 21665 96637 21711 96683
rect 21789 96637 21835 96683
rect 21913 96637 21959 96683
rect 22037 96637 22083 96683
rect 22161 96637 22207 96683
rect 22285 96637 22331 96683
rect 22409 96637 22455 96683
rect 22533 96637 22579 96683
rect 22657 96637 22703 96683
rect 22781 96637 22827 96683
rect 22905 96637 22951 96683
rect 23029 96637 23075 96683
rect 23153 96637 23199 96683
rect 23277 96637 23323 96683
rect 23401 96637 23447 96683
rect 23525 96637 23571 96683
rect 23649 96637 23695 96683
rect 23773 96637 23819 96683
rect 23897 96637 23943 96683
rect 24021 96637 24067 96683
rect 24145 96637 24191 96683
rect 24269 96637 24315 96683
rect 24393 96637 24439 96683
rect 24517 96637 24563 96683
rect 24641 96637 24687 96683
rect 24765 96637 24811 96683
rect 24889 96637 24935 96683
rect 25013 96637 25059 96683
rect 25137 96637 25183 96683
rect 25261 96637 25307 96683
rect 25385 96637 25431 96683
rect 25509 96637 25555 96683
rect 25633 96637 25679 96683
rect 25757 96637 25803 96683
rect 25881 96637 25927 96683
rect 26005 96637 26051 96683
rect 26129 96637 26175 96683
rect 26253 96637 26299 96683
rect 26377 96637 26423 96683
rect 26501 96637 26547 96683
rect 26625 96637 26671 96683
rect 26749 96637 26795 96683
rect 26873 96637 26919 96683
rect 26997 96637 27043 96683
rect 27121 96637 27167 96683
rect 27245 96637 27291 96683
rect 27369 96637 27415 96683
rect 27493 96637 27539 96683
rect 27617 96637 27663 96683
rect 27741 96637 27787 96683
rect 27865 96637 27911 96683
rect 27989 96637 28035 96683
rect 28113 96637 28159 96683
rect 28237 96637 28283 96683
rect 28361 96637 28407 96683
rect 28485 96637 28531 96683
rect 28609 96637 28655 96683
rect 28733 96637 28779 96683
rect 28857 96637 28903 96683
rect 28981 96637 29027 96683
rect 29105 96637 29151 96683
rect 29229 96637 29275 96683
rect 29353 96637 29399 96683
rect 29477 96637 29523 96683
rect 29601 96637 29647 96683
rect 29725 96637 29771 96683
rect 29849 96637 29895 96683
rect 29973 96637 30019 96683
rect 30097 96637 30143 96683
rect 30221 96637 30267 96683
rect 30345 96637 30391 96683
rect 30469 96637 30515 96683
rect 30593 96637 30639 96683
rect 30717 96637 30763 96683
rect 30841 96637 30887 96683
rect 30965 96637 31011 96683
rect 31089 96637 31135 96683
rect 31213 96637 31259 96683
rect 31337 96637 31383 96683
rect 31461 96637 31507 96683
rect 31585 96637 31631 96683
rect 31709 96637 31755 96683
rect 31833 96637 31879 96683
rect 31957 96637 32003 96683
rect 32081 96637 32127 96683
rect 32205 96637 32251 96683
rect 32329 96637 32375 96683
rect 32453 96637 32499 96683
rect 32577 96637 32623 96683
rect 32701 96637 32747 96683
rect 32825 96637 32871 96683
rect 32949 96637 32995 96683
rect 33073 96637 33119 96683
rect 33197 96637 33243 96683
rect 33321 96637 33367 96683
rect 33445 96637 33491 96683
rect 33569 96637 33615 96683
rect 33693 96637 33739 96683
rect 33817 96637 33863 96683
rect 33941 96637 33987 96683
rect 34065 96637 34111 96683
rect 34189 96637 34235 96683
rect 34313 96637 34359 96683
rect 34437 96637 34483 96683
rect 34561 96637 34607 96683
rect 34685 96637 34731 96683
rect 34809 96637 34855 96683
rect 34933 96637 34979 96683
rect 35057 96637 35103 96683
rect 35181 96637 35227 96683
rect 35305 96637 35351 96683
rect 35429 96637 35475 96683
rect 35553 96637 35599 96683
rect 35677 96637 35723 96683
rect 35801 96637 35847 96683
rect 35925 96637 35971 96683
rect 36049 96637 36095 96683
rect 36173 96637 36219 96683
rect 36297 96637 36343 96683
rect 36421 96637 36467 96683
rect 36545 96637 36591 96683
rect 36669 96637 36715 96683
rect 36793 96637 36839 96683
rect 36917 96637 36963 96683
rect 37041 96637 37087 96683
rect 37165 96637 37211 96683
rect 37289 96637 37335 96683
rect 37413 96637 37459 96683
rect 37537 96637 37583 96683
rect 37661 96637 37707 96683
rect 37785 96637 37831 96683
rect 37909 96637 37955 96683
rect 38033 96637 38079 96683
rect 38157 96637 38203 96683
rect 38281 96637 38327 96683
rect 38405 96637 38451 96683
rect 38529 96637 38575 96683
rect 38653 96637 38699 96683
rect 38777 96637 38823 96683
rect 38901 96637 38947 96683
rect 39025 96637 39071 96683
rect 39149 96637 39195 96683
rect 39273 96637 39319 96683
rect 39397 96637 39443 96683
rect 39521 96637 39567 96683
rect 39645 96637 39691 96683
rect 39769 96637 39815 96683
rect 39893 96637 39939 96683
rect 40017 96637 40063 96683
rect 40141 96637 40187 96683
rect 40265 96637 40311 96683
rect 40389 96637 40435 96683
rect 40513 96637 40559 96683
rect 40637 96637 40683 96683
rect 40761 96637 40807 96683
rect 40885 96637 40931 96683
rect 41009 96637 41055 96683
rect 41133 96637 41179 96683
rect 41257 96637 41303 96683
rect 41381 96637 41427 96683
rect 41505 96637 41551 96683
rect 41629 96637 41675 96683
rect 41753 96637 41799 96683
rect 41877 96637 41923 96683
rect 42001 96637 42047 96683
rect 42125 96637 42171 96683
rect 42249 96637 42295 96683
rect 42373 96637 42419 96683
rect 42497 96637 42543 96683
rect 42621 96637 42667 96683
rect 42745 96637 42791 96683
rect 42869 96637 42915 96683
rect 42993 96637 43039 96683
rect 43117 96637 43163 96683
rect 43241 96637 43287 96683
rect 43365 96637 43411 96683
rect 43489 96637 43535 96683
rect 43613 96637 43659 96683
rect 43737 96637 43783 96683
rect 43861 96637 43907 96683
rect 43985 96637 44031 96683
rect 44109 96637 44155 96683
rect 44233 96637 44279 96683
rect 44357 96637 44403 96683
rect 44481 96637 44527 96683
rect 44605 96637 44651 96683
rect 44729 96637 44775 96683
rect 44853 96637 44899 96683
rect 44977 96637 45023 96683
rect 45101 96637 45147 96683
rect 45225 96637 45271 96683
rect 45349 96637 45395 96683
rect 45473 96637 45519 96683
rect 45597 96637 45643 96683
rect 45721 96637 45767 96683
rect 45845 96637 45891 96683
rect 45969 96637 46015 96683
rect 46093 96637 46139 96683
rect 46217 96637 46263 96683
rect 46341 96637 46387 96683
rect 46465 96637 46511 96683
rect 46589 96637 46635 96683
rect 46713 96637 46759 96683
rect 46837 96637 46883 96683
rect 46961 96637 47007 96683
rect 47085 96637 47131 96683
rect 47209 96637 47255 96683
rect 47333 96637 47379 96683
rect 47457 96637 47503 96683
rect 47581 96637 47627 96683
rect 47705 96637 47751 96683
rect 47829 96637 47875 96683
rect 47953 96637 47999 96683
rect 48077 96637 48123 96683
rect 48201 96637 48247 96683
rect 48325 96637 48371 96683
rect 48449 96637 48495 96683
rect 48573 96637 48619 96683
rect 48697 96637 48743 96683
rect 48821 96637 48867 96683
rect 48945 96637 48991 96683
rect 49069 96637 49115 96683
rect 49193 96637 49239 96683
rect 49317 96637 49363 96683
rect 49441 96637 49487 96683
rect 49565 96637 49611 96683
rect 49689 96637 49735 96683
rect 49813 96637 49859 96683
rect 49937 96637 49983 96683
rect 50061 96637 50107 96683
rect 50185 96637 50231 96683
rect 50309 96637 50355 96683
rect 50433 96637 50479 96683
rect 50557 96637 50603 96683
rect 50681 96637 50727 96683
rect 50805 96637 50851 96683
rect 50929 96637 50975 96683
rect 51053 96637 51099 96683
rect 51177 96637 51223 96683
rect 51301 96637 51347 96683
rect 51425 96637 51471 96683
rect 51549 96637 51595 96683
rect 51673 96637 51719 96683
rect 51797 96637 51843 96683
rect 51921 96637 51967 96683
rect 52045 96637 52091 96683
rect 52169 96637 52215 96683
rect 52293 96637 52339 96683
rect 52417 96637 52463 96683
rect 52541 96637 52587 96683
rect 52665 96637 52711 96683
rect 52789 96637 52835 96683
rect 52913 96637 52959 96683
rect 53037 96637 53083 96683
rect 53161 96637 53207 96683
rect 53285 96637 53331 96683
rect 53409 96637 53455 96683
rect 53533 96637 53579 96683
rect 53657 96637 53703 96683
rect 53781 96637 53827 96683
rect 53905 96637 53951 96683
rect 54029 96637 54075 96683
rect 54153 96637 54199 96683
rect 54277 96637 54323 96683
rect 54401 96637 54447 96683
rect 54525 96637 54571 96683
rect 54649 96637 54695 96683
rect 54773 96637 54819 96683
rect 54897 96637 54943 96683
rect 55021 96637 55067 96683
rect 55145 96637 55191 96683
rect 55269 96637 55315 96683
rect 55393 96637 55439 96683
rect 55517 96637 55563 96683
rect 55641 96637 55687 96683
rect 55765 96637 55811 96683
rect 55889 96637 55935 96683
rect 56013 96637 56059 96683
rect 56137 96637 56183 96683
rect 56261 96637 56307 96683
rect 56385 96637 56431 96683
rect 56509 96637 56555 96683
rect 56633 96637 56679 96683
rect 56757 96637 56803 96683
rect 56881 96637 56927 96683
rect 57005 96637 57051 96683
rect 57129 96637 57175 96683
rect 57253 96637 57299 96683
rect 57377 96637 57423 96683
rect 57501 96637 57547 96683
rect 57625 96637 57671 96683
rect 57749 96637 57795 96683
rect 57873 96637 57919 96683
rect 57997 96637 58043 96683
rect 58121 96637 58167 96683
rect 58245 96637 58291 96683
rect 58369 96637 58415 96683
rect 58493 96637 58539 96683
rect 58617 96637 58663 96683
rect 58741 96637 58787 96683
rect 58865 96637 58911 96683
rect 58989 96637 59035 96683
rect 59113 96637 59159 96683
rect 59237 96637 59283 96683
rect 59361 96637 59407 96683
rect 59485 96637 59531 96683
rect 59609 96637 59655 96683
rect 59733 96637 59779 96683
rect 59857 96637 59903 96683
rect 59981 96637 60027 96683
rect 60105 96637 60151 96683
rect 60229 96637 60275 96683
rect 60353 96637 60399 96683
rect 60477 96637 60523 96683
rect 60601 96637 60647 96683
rect 60725 96637 60771 96683
rect 60849 96637 60895 96683
rect 60973 96637 61019 96683
rect 61097 96637 61143 96683
rect 61221 96637 61267 96683
rect 61345 96637 61391 96683
rect 61469 96637 61515 96683
rect 61593 96637 61639 96683
rect 61717 96637 61763 96683
rect 61841 96637 61887 96683
rect 61965 96637 62011 96683
rect 62089 96637 62135 96683
rect 62213 96637 62259 96683
rect 62337 96637 62383 96683
rect 62461 96637 62507 96683
rect 62585 96637 62631 96683
rect 62709 96637 62755 96683
rect 62833 96637 62879 96683
rect 62957 96637 63003 96683
rect 63081 96637 63127 96683
rect 63205 96637 63251 96683
rect 63329 96637 63375 96683
rect 63453 96637 63499 96683
rect 63577 96637 63623 96683
rect 63701 96637 63747 96683
rect 63825 96637 63871 96683
rect 63949 96637 63995 96683
rect 64073 96637 64119 96683
rect 64197 96637 64243 96683
rect 64321 96637 64367 96683
rect 64445 96637 64491 96683
rect 64569 96637 64615 96683
rect 64693 96637 64739 96683
rect 64817 96637 64863 96683
rect 64941 96637 64987 96683
rect 65065 96637 65111 96683
rect 65189 96637 65235 96683
rect 65313 96637 65359 96683
rect 65437 96637 65483 96683
rect 65561 96637 65607 96683
rect 65685 96637 65731 96683
rect 65809 96637 65855 96683
rect 65933 96637 65979 96683
rect 66057 96637 66103 96683
rect 66181 96637 66227 96683
rect 66305 96637 66351 96683
rect 66429 96637 66475 96683
rect 66553 96637 66599 96683
rect 66677 96637 66723 96683
rect 66801 96637 66847 96683
rect 66925 96637 66971 96683
rect 67049 96637 67095 96683
rect 67173 96637 67219 96683
rect 67297 96637 67343 96683
rect 67421 96637 67467 96683
rect 67545 96637 67591 96683
rect 67669 96637 67715 96683
rect 67793 96637 67839 96683
rect 67917 96637 67963 96683
rect 68041 96637 68087 96683
rect 68165 96637 68211 96683
rect 68289 96637 68335 96683
rect 68413 96637 68459 96683
rect 68537 96637 68583 96683
rect 68661 96637 68707 96683
rect 68785 96637 68831 96683
rect 68909 96637 68955 96683
rect 69033 96637 69079 96683
rect 69157 96637 69203 96683
rect 69281 96637 69327 96683
rect 69405 96637 69451 96683
rect 69529 96637 69575 96683
rect 69653 96637 69699 96683
rect 69777 96637 69823 96683
rect 69901 96637 69947 96683
rect 70025 96637 70071 96683
rect 70149 96637 70195 96683
rect 70273 96637 70319 96683
rect 70397 96637 70443 96683
rect 70521 96637 70567 96683
rect 70645 96637 70691 96683
rect 70769 96637 70815 96683
rect 70893 96637 70939 96683
rect 71017 96637 71063 96683
rect 71141 96637 71187 96683
rect 71265 96637 71311 96683
rect 71389 96637 71435 96683
rect 71513 96637 71559 96683
rect 71637 96637 71683 96683
rect 71761 96637 71807 96683
rect 71885 96637 71931 96683
rect 72009 96637 72055 96683
rect 72133 96637 72179 96683
rect 72257 96637 72303 96683
rect 72381 96637 72427 96683
rect 72505 96637 72551 96683
rect 72629 96637 72675 96683
rect 72753 96637 72799 96683
rect 72877 96637 72923 96683
rect 73001 96637 73047 96683
rect 73125 96637 73171 96683
rect 73249 96637 73295 96683
rect 73373 96637 73419 96683
rect 73497 96637 73543 96683
rect 73621 96637 73667 96683
rect 73745 96637 73791 96683
rect 73869 96637 73915 96683
rect 73993 96637 74039 96683
rect 74117 96637 74163 96683
rect 74241 96637 74287 96683
rect 74365 96637 74411 96683
rect 74489 96637 74535 96683
rect 74613 96637 74659 96683
rect 74737 96637 74783 96683
rect 74861 96637 74907 96683
rect 74985 96637 75031 96683
rect 75109 96637 75155 96683
rect 75233 96637 75279 96683
rect 75357 96637 75403 96683
rect 75481 96637 75527 96683
rect 75605 96637 75651 96683
rect 75729 96637 75775 96683
rect 75853 96637 75899 96683
rect 75977 96637 76023 96683
rect 76101 96637 76147 96683
rect 76225 96637 76271 96683
rect 76349 96637 76395 96683
rect 76473 96637 76519 96683
rect 76597 96637 76643 96683
rect 76721 96637 76767 96683
rect 76845 96637 76891 96683
rect 76969 96637 77015 96683
rect 77093 96637 77139 96683
rect 77217 96637 77263 96683
rect 77341 96637 77387 96683
rect 77465 96637 77511 96683
rect 77589 96637 77635 96683
rect 77713 96637 77759 96683
rect 77837 96637 77883 96683
rect 77961 96637 78007 96683
rect 78085 96637 78131 96683
rect 78209 96637 78255 96683
rect 78333 96637 78379 96683
rect 78457 96637 78503 96683
rect 78581 96637 78627 96683
rect 78705 96637 78751 96683
rect 78829 96637 78875 96683
rect 78953 96637 78999 96683
rect 79077 96637 79123 96683
rect 79201 96637 79247 96683
rect 79325 96637 79371 96683
rect 79449 96637 79495 96683
rect 79573 96637 79619 96683
rect 79697 96637 79743 96683
rect 79821 96637 79867 96683
rect 79945 96637 79991 96683
rect 80069 96637 80115 96683
rect 80193 96637 80239 96683
rect 80317 96637 80363 96683
rect 80441 96637 80487 96683
rect 80565 96637 80611 96683
rect 80689 96637 80735 96683
rect 80813 96637 80859 96683
rect 80937 96637 80983 96683
rect 81061 96637 81107 96683
rect 81185 96637 81231 96683
rect 81309 96637 81355 96683
rect 81433 96637 81479 96683
rect 81557 96637 81603 96683
rect 81681 96637 81727 96683
rect 81805 96637 81851 96683
rect 81929 96637 81975 96683
rect 82053 96637 82099 96683
rect 82177 96637 82223 96683
rect 82301 96637 82347 96683
rect 82425 96637 82471 96683
rect 82549 96637 82595 96683
rect 82673 96637 82719 96683
rect 82797 96637 82843 96683
rect 82921 96637 82967 96683
rect 83045 96637 83091 96683
rect 83169 96637 83215 96683
rect 83293 96637 83339 96683
rect 83417 96637 83463 96683
rect 83541 96637 83587 96683
rect 83665 96637 83711 96683
rect 83789 96637 83835 96683
rect 83913 96637 83959 96683
rect 84037 96637 84083 96683
rect 84161 96637 84207 96683
rect 84285 96637 84331 96683
rect 84409 96637 84455 96683
rect 84533 96637 84579 96683
rect 84657 96637 84703 96683
rect 84781 96637 84827 96683
rect 84905 96637 84951 96683
rect 85029 96637 85075 96683
rect 85153 96637 85199 96683
rect 85277 96637 85323 96683
rect 85401 96637 85447 96683
rect 85525 96637 85571 96683
rect 85649 96637 85695 96683
rect 89 96513 135 96559
rect 213 96513 259 96559
rect 337 96513 383 96559
rect 461 96513 507 96559
rect 585 96513 631 96559
rect 709 96513 755 96559
rect 833 96513 879 96559
rect 957 96513 1003 96559
rect 1081 96513 1127 96559
rect 1205 96513 1251 96559
rect 1329 96513 1375 96559
rect 1453 96513 1499 96559
rect 1577 96513 1623 96559
rect 1701 96513 1747 96559
rect 1825 96513 1871 96559
rect 1949 96513 1995 96559
rect 2073 96513 2119 96559
rect 2197 96513 2243 96559
rect 2321 96513 2367 96559
rect 2445 96513 2491 96559
rect 2569 96513 2615 96559
rect 2693 96513 2739 96559
rect 2817 96513 2863 96559
rect 2941 96513 2987 96559
rect 3065 96513 3111 96559
rect 3189 96513 3235 96559
rect 3313 96513 3359 96559
rect 3437 96513 3483 96559
rect 3561 96513 3607 96559
rect 3685 96513 3731 96559
rect 3809 96513 3855 96559
rect 3933 96513 3979 96559
rect 4057 96513 4103 96559
rect 4181 96513 4227 96559
rect 4305 96513 4351 96559
rect 4429 96513 4475 96559
rect 4553 96513 4599 96559
rect 4677 96513 4723 96559
rect 4801 96513 4847 96559
rect 4925 96513 4971 96559
rect 5049 96513 5095 96559
rect 5173 96513 5219 96559
rect 5297 96513 5343 96559
rect 5421 96513 5467 96559
rect 5545 96513 5591 96559
rect 5669 96513 5715 96559
rect 5793 96513 5839 96559
rect 5917 96513 5963 96559
rect 6041 96513 6087 96559
rect 6165 96513 6211 96559
rect 6289 96513 6335 96559
rect 6413 96513 6459 96559
rect 6537 96513 6583 96559
rect 6661 96513 6707 96559
rect 6785 96513 6831 96559
rect 6909 96513 6955 96559
rect 7033 96513 7079 96559
rect 7157 96513 7203 96559
rect 7281 96513 7327 96559
rect 7405 96513 7451 96559
rect 7529 96513 7575 96559
rect 7653 96513 7699 96559
rect 7777 96513 7823 96559
rect 7901 96513 7947 96559
rect 8025 96513 8071 96559
rect 8149 96513 8195 96559
rect 8273 96513 8319 96559
rect 8397 96513 8443 96559
rect 8521 96513 8567 96559
rect 8645 96513 8691 96559
rect 8769 96513 8815 96559
rect 8893 96513 8939 96559
rect 9017 96513 9063 96559
rect 9141 96513 9187 96559
rect 9265 96513 9311 96559
rect 9389 96513 9435 96559
rect 9513 96513 9559 96559
rect 9637 96513 9683 96559
rect 9761 96513 9807 96559
rect 9885 96513 9931 96559
rect 10009 96513 10055 96559
rect 10133 96513 10179 96559
rect 10257 96513 10303 96559
rect 10381 96513 10427 96559
rect 10505 96513 10551 96559
rect 10629 96513 10675 96559
rect 10753 96513 10799 96559
rect 10877 96513 10923 96559
rect 11001 96513 11047 96559
rect 11125 96513 11171 96559
rect 11249 96513 11295 96559
rect 11373 96513 11419 96559
rect 11497 96513 11543 96559
rect 11621 96513 11667 96559
rect 11745 96513 11791 96559
rect 11869 96513 11915 96559
rect 11993 96513 12039 96559
rect 12117 96513 12163 96559
rect 12241 96513 12287 96559
rect 12365 96513 12411 96559
rect 12489 96513 12535 96559
rect 12613 96513 12659 96559
rect 12737 96513 12783 96559
rect 12861 96513 12907 96559
rect 12985 96513 13031 96559
rect 13109 96513 13155 96559
rect 13233 96513 13279 96559
rect 13357 96513 13403 96559
rect 13481 96513 13527 96559
rect 13605 96513 13651 96559
rect 13729 96513 13775 96559
rect 13853 96513 13899 96559
rect 13977 96513 14023 96559
rect 14101 96513 14147 96559
rect 14225 96513 14271 96559
rect 14349 96513 14395 96559
rect 14473 96513 14519 96559
rect 14597 96513 14643 96559
rect 14721 96513 14767 96559
rect 14845 96513 14891 96559
rect 14969 96513 15015 96559
rect 15093 96513 15139 96559
rect 15217 96513 15263 96559
rect 15341 96513 15387 96559
rect 15465 96513 15511 96559
rect 15589 96513 15635 96559
rect 15713 96513 15759 96559
rect 15837 96513 15883 96559
rect 15961 96513 16007 96559
rect 16085 96513 16131 96559
rect 16209 96513 16255 96559
rect 16333 96513 16379 96559
rect 16457 96513 16503 96559
rect 16581 96513 16627 96559
rect 16705 96513 16751 96559
rect 16829 96513 16875 96559
rect 16953 96513 16999 96559
rect 17077 96513 17123 96559
rect 17201 96513 17247 96559
rect 17325 96513 17371 96559
rect 17449 96513 17495 96559
rect 17573 96513 17619 96559
rect 17697 96513 17743 96559
rect 17821 96513 17867 96559
rect 17945 96513 17991 96559
rect 18069 96513 18115 96559
rect 18193 96513 18239 96559
rect 18317 96513 18363 96559
rect 18441 96513 18487 96559
rect 18565 96513 18611 96559
rect 18689 96513 18735 96559
rect 18813 96513 18859 96559
rect 18937 96513 18983 96559
rect 19061 96513 19107 96559
rect 19185 96513 19231 96559
rect 19309 96513 19355 96559
rect 19433 96513 19479 96559
rect 19557 96513 19603 96559
rect 19681 96513 19727 96559
rect 19805 96513 19851 96559
rect 19929 96513 19975 96559
rect 20053 96513 20099 96559
rect 20177 96513 20223 96559
rect 20301 96513 20347 96559
rect 20425 96513 20471 96559
rect 20549 96513 20595 96559
rect 20673 96513 20719 96559
rect 20797 96513 20843 96559
rect 20921 96513 20967 96559
rect 21045 96513 21091 96559
rect 21169 96513 21215 96559
rect 21293 96513 21339 96559
rect 21417 96513 21463 96559
rect 21541 96513 21587 96559
rect 21665 96513 21711 96559
rect 21789 96513 21835 96559
rect 21913 96513 21959 96559
rect 22037 96513 22083 96559
rect 22161 96513 22207 96559
rect 22285 96513 22331 96559
rect 22409 96513 22455 96559
rect 22533 96513 22579 96559
rect 22657 96513 22703 96559
rect 22781 96513 22827 96559
rect 22905 96513 22951 96559
rect 23029 96513 23075 96559
rect 23153 96513 23199 96559
rect 23277 96513 23323 96559
rect 23401 96513 23447 96559
rect 23525 96513 23571 96559
rect 23649 96513 23695 96559
rect 23773 96513 23819 96559
rect 23897 96513 23943 96559
rect 24021 96513 24067 96559
rect 24145 96513 24191 96559
rect 24269 96513 24315 96559
rect 24393 96513 24439 96559
rect 24517 96513 24563 96559
rect 24641 96513 24687 96559
rect 24765 96513 24811 96559
rect 24889 96513 24935 96559
rect 25013 96513 25059 96559
rect 25137 96513 25183 96559
rect 25261 96513 25307 96559
rect 25385 96513 25431 96559
rect 25509 96513 25555 96559
rect 25633 96513 25679 96559
rect 25757 96513 25803 96559
rect 25881 96513 25927 96559
rect 26005 96513 26051 96559
rect 26129 96513 26175 96559
rect 26253 96513 26299 96559
rect 26377 96513 26423 96559
rect 26501 96513 26547 96559
rect 26625 96513 26671 96559
rect 26749 96513 26795 96559
rect 26873 96513 26919 96559
rect 26997 96513 27043 96559
rect 27121 96513 27167 96559
rect 27245 96513 27291 96559
rect 27369 96513 27415 96559
rect 27493 96513 27539 96559
rect 27617 96513 27663 96559
rect 27741 96513 27787 96559
rect 27865 96513 27911 96559
rect 27989 96513 28035 96559
rect 28113 96513 28159 96559
rect 28237 96513 28283 96559
rect 28361 96513 28407 96559
rect 28485 96513 28531 96559
rect 28609 96513 28655 96559
rect 28733 96513 28779 96559
rect 28857 96513 28903 96559
rect 28981 96513 29027 96559
rect 29105 96513 29151 96559
rect 29229 96513 29275 96559
rect 29353 96513 29399 96559
rect 29477 96513 29523 96559
rect 29601 96513 29647 96559
rect 29725 96513 29771 96559
rect 29849 96513 29895 96559
rect 29973 96513 30019 96559
rect 30097 96513 30143 96559
rect 30221 96513 30267 96559
rect 30345 96513 30391 96559
rect 30469 96513 30515 96559
rect 30593 96513 30639 96559
rect 30717 96513 30763 96559
rect 30841 96513 30887 96559
rect 30965 96513 31011 96559
rect 31089 96513 31135 96559
rect 31213 96513 31259 96559
rect 31337 96513 31383 96559
rect 31461 96513 31507 96559
rect 31585 96513 31631 96559
rect 31709 96513 31755 96559
rect 31833 96513 31879 96559
rect 31957 96513 32003 96559
rect 32081 96513 32127 96559
rect 32205 96513 32251 96559
rect 32329 96513 32375 96559
rect 32453 96513 32499 96559
rect 32577 96513 32623 96559
rect 32701 96513 32747 96559
rect 32825 96513 32871 96559
rect 32949 96513 32995 96559
rect 33073 96513 33119 96559
rect 33197 96513 33243 96559
rect 33321 96513 33367 96559
rect 33445 96513 33491 96559
rect 33569 96513 33615 96559
rect 33693 96513 33739 96559
rect 33817 96513 33863 96559
rect 33941 96513 33987 96559
rect 34065 96513 34111 96559
rect 34189 96513 34235 96559
rect 34313 96513 34359 96559
rect 34437 96513 34483 96559
rect 34561 96513 34607 96559
rect 34685 96513 34731 96559
rect 34809 96513 34855 96559
rect 34933 96513 34979 96559
rect 35057 96513 35103 96559
rect 35181 96513 35227 96559
rect 35305 96513 35351 96559
rect 35429 96513 35475 96559
rect 35553 96513 35599 96559
rect 35677 96513 35723 96559
rect 35801 96513 35847 96559
rect 35925 96513 35971 96559
rect 36049 96513 36095 96559
rect 36173 96513 36219 96559
rect 36297 96513 36343 96559
rect 36421 96513 36467 96559
rect 36545 96513 36591 96559
rect 36669 96513 36715 96559
rect 36793 96513 36839 96559
rect 36917 96513 36963 96559
rect 37041 96513 37087 96559
rect 37165 96513 37211 96559
rect 37289 96513 37335 96559
rect 37413 96513 37459 96559
rect 37537 96513 37583 96559
rect 37661 96513 37707 96559
rect 37785 96513 37831 96559
rect 37909 96513 37955 96559
rect 38033 96513 38079 96559
rect 38157 96513 38203 96559
rect 38281 96513 38327 96559
rect 38405 96513 38451 96559
rect 38529 96513 38575 96559
rect 38653 96513 38699 96559
rect 38777 96513 38823 96559
rect 38901 96513 38947 96559
rect 39025 96513 39071 96559
rect 39149 96513 39195 96559
rect 39273 96513 39319 96559
rect 39397 96513 39443 96559
rect 39521 96513 39567 96559
rect 39645 96513 39691 96559
rect 39769 96513 39815 96559
rect 39893 96513 39939 96559
rect 40017 96513 40063 96559
rect 40141 96513 40187 96559
rect 40265 96513 40311 96559
rect 40389 96513 40435 96559
rect 40513 96513 40559 96559
rect 40637 96513 40683 96559
rect 40761 96513 40807 96559
rect 40885 96513 40931 96559
rect 41009 96513 41055 96559
rect 41133 96513 41179 96559
rect 41257 96513 41303 96559
rect 41381 96513 41427 96559
rect 41505 96513 41551 96559
rect 41629 96513 41675 96559
rect 41753 96513 41799 96559
rect 41877 96513 41923 96559
rect 42001 96513 42047 96559
rect 42125 96513 42171 96559
rect 42249 96513 42295 96559
rect 42373 96513 42419 96559
rect 42497 96513 42543 96559
rect 42621 96513 42667 96559
rect 42745 96513 42791 96559
rect 42869 96513 42915 96559
rect 42993 96513 43039 96559
rect 43117 96513 43163 96559
rect 43241 96513 43287 96559
rect 43365 96513 43411 96559
rect 43489 96513 43535 96559
rect 43613 96513 43659 96559
rect 43737 96513 43783 96559
rect 43861 96513 43907 96559
rect 43985 96513 44031 96559
rect 44109 96513 44155 96559
rect 44233 96513 44279 96559
rect 44357 96513 44403 96559
rect 44481 96513 44527 96559
rect 44605 96513 44651 96559
rect 44729 96513 44775 96559
rect 44853 96513 44899 96559
rect 44977 96513 45023 96559
rect 45101 96513 45147 96559
rect 45225 96513 45271 96559
rect 45349 96513 45395 96559
rect 45473 96513 45519 96559
rect 45597 96513 45643 96559
rect 45721 96513 45767 96559
rect 45845 96513 45891 96559
rect 45969 96513 46015 96559
rect 46093 96513 46139 96559
rect 46217 96513 46263 96559
rect 46341 96513 46387 96559
rect 46465 96513 46511 96559
rect 46589 96513 46635 96559
rect 46713 96513 46759 96559
rect 46837 96513 46883 96559
rect 46961 96513 47007 96559
rect 47085 96513 47131 96559
rect 47209 96513 47255 96559
rect 47333 96513 47379 96559
rect 47457 96513 47503 96559
rect 47581 96513 47627 96559
rect 47705 96513 47751 96559
rect 47829 96513 47875 96559
rect 47953 96513 47999 96559
rect 48077 96513 48123 96559
rect 48201 96513 48247 96559
rect 48325 96513 48371 96559
rect 48449 96513 48495 96559
rect 48573 96513 48619 96559
rect 48697 96513 48743 96559
rect 48821 96513 48867 96559
rect 48945 96513 48991 96559
rect 49069 96513 49115 96559
rect 49193 96513 49239 96559
rect 49317 96513 49363 96559
rect 49441 96513 49487 96559
rect 49565 96513 49611 96559
rect 49689 96513 49735 96559
rect 49813 96513 49859 96559
rect 49937 96513 49983 96559
rect 50061 96513 50107 96559
rect 50185 96513 50231 96559
rect 50309 96513 50355 96559
rect 50433 96513 50479 96559
rect 50557 96513 50603 96559
rect 50681 96513 50727 96559
rect 50805 96513 50851 96559
rect 50929 96513 50975 96559
rect 51053 96513 51099 96559
rect 51177 96513 51223 96559
rect 51301 96513 51347 96559
rect 51425 96513 51471 96559
rect 51549 96513 51595 96559
rect 51673 96513 51719 96559
rect 51797 96513 51843 96559
rect 51921 96513 51967 96559
rect 52045 96513 52091 96559
rect 52169 96513 52215 96559
rect 52293 96513 52339 96559
rect 52417 96513 52463 96559
rect 52541 96513 52587 96559
rect 52665 96513 52711 96559
rect 52789 96513 52835 96559
rect 52913 96513 52959 96559
rect 53037 96513 53083 96559
rect 53161 96513 53207 96559
rect 53285 96513 53331 96559
rect 53409 96513 53455 96559
rect 53533 96513 53579 96559
rect 53657 96513 53703 96559
rect 53781 96513 53827 96559
rect 53905 96513 53951 96559
rect 54029 96513 54075 96559
rect 54153 96513 54199 96559
rect 54277 96513 54323 96559
rect 54401 96513 54447 96559
rect 54525 96513 54571 96559
rect 54649 96513 54695 96559
rect 54773 96513 54819 96559
rect 54897 96513 54943 96559
rect 55021 96513 55067 96559
rect 55145 96513 55191 96559
rect 55269 96513 55315 96559
rect 55393 96513 55439 96559
rect 55517 96513 55563 96559
rect 55641 96513 55687 96559
rect 55765 96513 55811 96559
rect 55889 96513 55935 96559
rect 56013 96513 56059 96559
rect 56137 96513 56183 96559
rect 56261 96513 56307 96559
rect 56385 96513 56431 96559
rect 56509 96513 56555 96559
rect 56633 96513 56679 96559
rect 56757 96513 56803 96559
rect 56881 96513 56927 96559
rect 57005 96513 57051 96559
rect 57129 96513 57175 96559
rect 57253 96513 57299 96559
rect 57377 96513 57423 96559
rect 57501 96513 57547 96559
rect 57625 96513 57671 96559
rect 57749 96513 57795 96559
rect 57873 96513 57919 96559
rect 57997 96513 58043 96559
rect 58121 96513 58167 96559
rect 58245 96513 58291 96559
rect 58369 96513 58415 96559
rect 58493 96513 58539 96559
rect 58617 96513 58663 96559
rect 58741 96513 58787 96559
rect 58865 96513 58911 96559
rect 58989 96513 59035 96559
rect 59113 96513 59159 96559
rect 59237 96513 59283 96559
rect 59361 96513 59407 96559
rect 59485 96513 59531 96559
rect 59609 96513 59655 96559
rect 59733 96513 59779 96559
rect 59857 96513 59903 96559
rect 59981 96513 60027 96559
rect 60105 96513 60151 96559
rect 60229 96513 60275 96559
rect 60353 96513 60399 96559
rect 60477 96513 60523 96559
rect 60601 96513 60647 96559
rect 60725 96513 60771 96559
rect 60849 96513 60895 96559
rect 60973 96513 61019 96559
rect 61097 96513 61143 96559
rect 61221 96513 61267 96559
rect 61345 96513 61391 96559
rect 61469 96513 61515 96559
rect 61593 96513 61639 96559
rect 61717 96513 61763 96559
rect 61841 96513 61887 96559
rect 61965 96513 62011 96559
rect 62089 96513 62135 96559
rect 62213 96513 62259 96559
rect 62337 96513 62383 96559
rect 62461 96513 62507 96559
rect 62585 96513 62631 96559
rect 62709 96513 62755 96559
rect 62833 96513 62879 96559
rect 62957 96513 63003 96559
rect 63081 96513 63127 96559
rect 63205 96513 63251 96559
rect 63329 96513 63375 96559
rect 63453 96513 63499 96559
rect 63577 96513 63623 96559
rect 63701 96513 63747 96559
rect 63825 96513 63871 96559
rect 63949 96513 63995 96559
rect 64073 96513 64119 96559
rect 64197 96513 64243 96559
rect 64321 96513 64367 96559
rect 64445 96513 64491 96559
rect 64569 96513 64615 96559
rect 64693 96513 64739 96559
rect 64817 96513 64863 96559
rect 64941 96513 64987 96559
rect 65065 96513 65111 96559
rect 65189 96513 65235 96559
rect 65313 96513 65359 96559
rect 65437 96513 65483 96559
rect 65561 96513 65607 96559
rect 65685 96513 65731 96559
rect 65809 96513 65855 96559
rect 65933 96513 65979 96559
rect 66057 96513 66103 96559
rect 66181 96513 66227 96559
rect 66305 96513 66351 96559
rect 66429 96513 66475 96559
rect 66553 96513 66599 96559
rect 66677 96513 66723 96559
rect 66801 96513 66847 96559
rect 66925 96513 66971 96559
rect 67049 96513 67095 96559
rect 67173 96513 67219 96559
rect 67297 96513 67343 96559
rect 67421 96513 67467 96559
rect 67545 96513 67591 96559
rect 67669 96513 67715 96559
rect 67793 96513 67839 96559
rect 67917 96513 67963 96559
rect 68041 96513 68087 96559
rect 68165 96513 68211 96559
rect 68289 96513 68335 96559
rect 68413 96513 68459 96559
rect 68537 96513 68583 96559
rect 68661 96513 68707 96559
rect 68785 96513 68831 96559
rect 68909 96513 68955 96559
rect 69033 96513 69079 96559
rect 69157 96513 69203 96559
rect 69281 96513 69327 96559
rect 69405 96513 69451 96559
rect 69529 96513 69575 96559
rect 69653 96513 69699 96559
rect 69777 96513 69823 96559
rect 69901 96513 69947 96559
rect 70025 96513 70071 96559
rect 70149 96513 70195 96559
rect 70273 96513 70319 96559
rect 70397 96513 70443 96559
rect 70521 96513 70567 96559
rect 70645 96513 70691 96559
rect 70769 96513 70815 96559
rect 70893 96513 70939 96559
rect 71017 96513 71063 96559
rect 71141 96513 71187 96559
rect 71265 96513 71311 96559
rect 71389 96513 71435 96559
rect 71513 96513 71559 96559
rect 71637 96513 71683 96559
rect 71761 96513 71807 96559
rect 71885 96513 71931 96559
rect 72009 96513 72055 96559
rect 72133 96513 72179 96559
rect 72257 96513 72303 96559
rect 72381 96513 72427 96559
rect 72505 96513 72551 96559
rect 72629 96513 72675 96559
rect 72753 96513 72799 96559
rect 72877 96513 72923 96559
rect 73001 96513 73047 96559
rect 73125 96513 73171 96559
rect 73249 96513 73295 96559
rect 73373 96513 73419 96559
rect 73497 96513 73543 96559
rect 73621 96513 73667 96559
rect 73745 96513 73791 96559
rect 73869 96513 73915 96559
rect 73993 96513 74039 96559
rect 74117 96513 74163 96559
rect 74241 96513 74287 96559
rect 74365 96513 74411 96559
rect 74489 96513 74535 96559
rect 74613 96513 74659 96559
rect 74737 96513 74783 96559
rect 74861 96513 74907 96559
rect 74985 96513 75031 96559
rect 75109 96513 75155 96559
rect 75233 96513 75279 96559
rect 75357 96513 75403 96559
rect 75481 96513 75527 96559
rect 75605 96513 75651 96559
rect 75729 96513 75775 96559
rect 75853 96513 75899 96559
rect 75977 96513 76023 96559
rect 76101 96513 76147 96559
rect 76225 96513 76271 96559
rect 76349 96513 76395 96559
rect 76473 96513 76519 96559
rect 76597 96513 76643 96559
rect 76721 96513 76767 96559
rect 76845 96513 76891 96559
rect 76969 96513 77015 96559
rect 77093 96513 77139 96559
rect 77217 96513 77263 96559
rect 77341 96513 77387 96559
rect 77465 96513 77511 96559
rect 77589 96513 77635 96559
rect 77713 96513 77759 96559
rect 77837 96513 77883 96559
rect 77961 96513 78007 96559
rect 78085 96513 78131 96559
rect 78209 96513 78255 96559
rect 78333 96513 78379 96559
rect 78457 96513 78503 96559
rect 78581 96513 78627 96559
rect 78705 96513 78751 96559
rect 78829 96513 78875 96559
rect 78953 96513 78999 96559
rect 79077 96513 79123 96559
rect 79201 96513 79247 96559
rect 79325 96513 79371 96559
rect 79449 96513 79495 96559
rect 79573 96513 79619 96559
rect 79697 96513 79743 96559
rect 79821 96513 79867 96559
rect 79945 96513 79991 96559
rect 80069 96513 80115 96559
rect 80193 96513 80239 96559
rect 80317 96513 80363 96559
rect 80441 96513 80487 96559
rect 80565 96513 80611 96559
rect 80689 96513 80735 96559
rect 80813 96513 80859 96559
rect 80937 96513 80983 96559
rect 81061 96513 81107 96559
rect 81185 96513 81231 96559
rect 81309 96513 81355 96559
rect 81433 96513 81479 96559
rect 81557 96513 81603 96559
rect 81681 96513 81727 96559
rect 81805 96513 81851 96559
rect 81929 96513 81975 96559
rect 82053 96513 82099 96559
rect 82177 96513 82223 96559
rect 82301 96513 82347 96559
rect 82425 96513 82471 96559
rect 82549 96513 82595 96559
rect 82673 96513 82719 96559
rect 82797 96513 82843 96559
rect 82921 96513 82967 96559
rect 83045 96513 83091 96559
rect 83169 96513 83215 96559
rect 83293 96513 83339 96559
rect 83417 96513 83463 96559
rect 83541 96513 83587 96559
rect 83665 96513 83711 96559
rect 83789 96513 83835 96559
rect 83913 96513 83959 96559
rect 84037 96513 84083 96559
rect 84161 96513 84207 96559
rect 84285 96513 84331 96559
rect 84409 96513 84455 96559
rect 84533 96513 84579 96559
rect 84657 96513 84703 96559
rect 84781 96513 84827 96559
rect 84905 96513 84951 96559
rect 85029 96513 85075 96559
rect 85153 96513 85199 96559
rect 85277 96513 85323 96559
rect 85401 96513 85447 96559
rect 85525 96513 85571 96559
rect 85649 96513 85695 96559
rect 89 96389 135 96435
rect 213 96389 259 96435
rect 337 96389 383 96435
rect 461 96389 507 96435
rect 585 96389 631 96435
rect 709 96389 755 96435
rect 833 96389 879 96435
rect 957 96389 1003 96435
rect 1081 96389 1127 96435
rect 1205 96389 1251 96435
rect 1329 96389 1375 96435
rect 1453 96389 1499 96435
rect 1577 96389 1623 96435
rect 1701 96389 1747 96435
rect 1825 96389 1871 96435
rect 1949 96389 1995 96435
rect 2073 96389 2119 96435
rect 2197 96389 2243 96435
rect 2321 96389 2367 96435
rect 2445 96389 2491 96435
rect 2569 96389 2615 96435
rect 2693 96389 2739 96435
rect 2817 96389 2863 96435
rect 2941 96389 2987 96435
rect 3065 96389 3111 96435
rect 3189 96389 3235 96435
rect 3313 96389 3359 96435
rect 3437 96389 3483 96435
rect 3561 96389 3607 96435
rect 3685 96389 3731 96435
rect 3809 96389 3855 96435
rect 3933 96389 3979 96435
rect 4057 96389 4103 96435
rect 4181 96389 4227 96435
rect 4305 96389 4351 96435
rect 4429 96389 4475 96435
rect 4553 96389 4599 96435
rect 4677 96389 4723 96435
rect 4801 96389 4847 96435
rect 4925 96389 4971 96435
rect 5049 96389 5095 96435
rect 5173 96389 5219 96435
rect 5297 96389 5343 96435
rect 5421 96389 5467 96435
rect 5545 96389 5591 96435
rect 5669 96389 5715 96435
rect 5793 96389 5839 96435
rect 5917 96389 5963 96435
rect 6041 96389 6087 96435
rect 6165 96389 6211 96435
rect 6289 96389 6335 96435
rect 6413 96389 6459 96435
rect 6537 96389 6583 96435
rect 6661 96389 6707 96435
rect 6785 96389 6831 96435
rect 6909 96389 6955 96435
rect 7033 96389 7079 96435
rect 7157 96389 7203 96435
rect 7281 96389 7327 96435
rect 7405 96389 7451 96435
rect 7529 96389 7575 96435
rect 7653 96389 7699 96435
rect 7777 96389 7823 96435
rect 7901 96389 7947 96435
rect 8025 96389 8071 96435
rect 8149 96389 8195 96435
rect 8273 96389 8319 96435
rect 8397 96389 8443 96435
rect 8521 96389 8567 96435
rect 8645 96389 8691 96435
rect 8769 96389 8815 96435
rect 8893 96389 8939 96435
rect 9017 96389 9063 96435
rect 9141 96389 9187 96435
rect 9265 96389 9311 96435
rect 9389 96389 9435 96435
rect 9513 96389 9559 96435
rect 9637 96389 9683 96435
rect 9761 96389 9807 96435
rect 9885 96389 9931 96435
rect 10009 96389 10055 96435
rect 10133 96389 10179 96435
rect 10257 96389 10303 96435
rect 10381 96389 10427 96435
rect 10505 96389 10551 96435
rect 10629 96389 10675 96435
rect 10753 96389 10799 96435
rect 10877 96389 10923 96435
rect 11001 96389 11047 96435
rect 11125 96389 11171 96435
rect 11249 96389 11295 96435
rect 11373 96389 11419 96435
rect 11497 96389 11543 96435
rect 11621 96389 11667 96435
rect 11745 96389 11791 96435
rect 11869 96389 11915 96435
rect 11993 96389 12039 96435
rect 12117 96389 12163 96435
rect 12241 96389 12287 96435
rect 12365 96389 12411 96435
rect 12489 96389 12535 96435
rect 12613 96389 12659 96435
rect 12737 96389 12783 96435
rect 12861 96389 12907 96435
rect 12985 96389 13031 96435
rect 13109 96389 13155 96435
rect 13233 96389 13279 96435
rect 13357 96389 13403 96435
rect 13481 96389 13527 96435
rect 13605 96389 13651 96435
rect 13729 96389 13775 96435
rect 13853 96389 13899 96435
rect 13977 96389 14023 96435
rect 14101 96389 14147 96435
rect 14225 96389 14271 96435
rect 14349 96389 14395 96435
rect 14473 96389 14519 96435
rect 14597 96389 14643 96435
rect 14721 96389 14767 96435
rect 14845 96389 14891 96435
rect 14969 96389 15015 96435
rect 15093 96389 15139 96435
rect 15217 96389 15263 96435
rect 15341 96389 15387 96435
rect 15465 96389 15511 96435
rect 15589 96389 15635 96435
rect 15713 96389 15759 96435
rect 15837 96389 15883 96435
rect 15961 96389 16007 96435
rect 16085 96389 16131 96435
rect 16209 96389 16255 96435
rect 16333 96389 16379 96435
rect 16457 96389 16503 96435
rect 16581 96389 16627 96435
rect 16705 96389 16751 96435
rect 16829 96389 16875 96435
rect 16953 96389 16999 96435
rect 17077 96389 17123 96435
rect 17201 96389 17247 96435
rect 17325 96389 17371 96435
rect 17449 96389 17495 96435
rect 17573 96389 17619 96435
rect 17697 96389 17743 96435
rect 17821 96389 17867 96435
rect 17945 96389 17991 96435
rect 18069 96389 18115 96435
rect 18193 96389 18239 96435
rect 18317 96389 18363 96435
rect 18441 96389 18487 96435
rect 18565 96389 18611 96435
rect 18689 96389 18735 96435
rect 18813 96389 18859 96435
rect 18937 96389 18983 96435
rect 19061 96389 19107 96435
rect 19185 96389 19231 96435
rect 19309 96389 19355 96435
rect 19433 96389 19479 96435
rect 19557 96389 19603 96435
rect 19681 96389 19727 96435
rect 19805 96389 19851 96435
rect 19929 96389 19975 96435
rect 20053 96389 20099 96435
rect 20177 96389 20223 96435
rect 20301 96389 20347 96435
rect 20425 96389 20471 96435
rect 20549 96389 20595 96435
rect 20673 96389 20719 96435
rect 20797 96389 20843 96435
rect 20921 96389 20967 96435
rect 21045 96389 21091 96435
rect 21169 96389 21215 96435
rect 21293 96389 21339 96435
rect 21417 96389 21463 96435
rect 21541 96389 21587 96435
rect 21665 96389 21711 96435
rect 21789 96389 21835 96435
rect 21913 96389 21959 96435
rect 22037 96389 22083 96435
rect 22161 96389 22207 96435
rect 22285 96389 22331 96435
rect 22409 96389 22455 96435
rect 22533 96389 22579 96435
rect 22657 96389 22703 96435
rect 22781 96389 22827 96435
rect 22905 96389 22951 96435
rect 23029 96389 23075 96435
rect 23153 96389 23199 96435
rect 23277 96389 23323 96435
rect 23401 96389 23447 96435
rect 23525 96389 23571 96435
rect 23649 96389 23695 96435
rect 23773 96389 23819 96435
rect 23897 96389 23943 96435
rect 24021 96389 24067 96435
rect 24145 96389 24191 96435
rect 24269 96389 24315 96435
rect 24393 96389 24439 96435
rect 24517 96389 24563 96435
rect 24641 96389 24687 96435
rect 24765 96389 24811 96435
rect 24889 96389 24935 96435
rect 25013 96389 25059 96435
rect 25137 96389 25183 96435
rect 25261 96389 25307 96435
rect 25385 96389 25431 96435
rect 25509 96389 25555 96435
rect 25633 96389 25679 96435
rect 25757 96389 25803 96435
rect 25881 96389 25927 96435
rect 26005 96389 26051 96435
rect 26129 96389 26175 96435
rect 26253 96389 26299 96435
rect 26377 96389 26423 96435
rect 26501 96389 26547 96435
rect 26625 96389 26671 96435
rect 26749 96389 26795 96435
rect 26873 96389 26919 96435
rect 26997 96389 27043 96435
rect 27121 96389 27167 96435
rect 27245 96389 27291 96435
rect 27369 96389 27415 96435
rect 27493 96389 27539 96435
rect 27617 96389 27663 96435
rect 27741 96389 27787 96435
rect 27865 96389 27911 96435
rect 27989 96389 28035 96435
rect 28113 96389 28159 96435
rect 28237 96389 28283 96435
rect 28361 96389 28407 96435
rect 28485 96389 28531 96435
rect 28609 96389 28655 96435
rect 28733 96389 28779 96435
rect 28857 96389 28903 96435
rect 28981 96389 29027 96435
rect 29105 96389 29151 96435
rect 29229 96389 29275 96435
rect 29353 96389 29399 96435
rect 29477 96389 29523 96435
rect 29601 96389 29647 96435
rect 29725 96389 29771 96435
rect 29849 96389 29895 96435
rect 29973 96389 30019 96435
rect 30097 96389 30143 96435
rect 30221 96389 30267 96435
rect 30345 96389 30391 96435
rect 30469 96389 30515 96435
rect 30593 96389 30639 96435
rect 30717 96389 30763 96435
rect 30841 96389 30887 96435
rect 30965 96389 31011 96435
rect 31089 96389 31135 96435
rect 31213 96389 31259 96435
rect 31337 96389 31383 96435
rect 31461 96389 31507 96435
rect 31585 96389 31631 96435
rect 31709 96389 31755 96435
rect 31833 96389 31879 96435
rect 31957 96389 32003 96435
rect 32081 96389 32127 96435
rect 32205 96389 32251 96435
rect 32329 96389 32375 96435
rect 32453 96389 32499 96435
rect 32577 96389 32623 96435
rect 32701 96389 32747 96435
rect 32825 96389 32871 96435
rect 32949 96389 32995 96435
rect 33073 96389 33119 96435
rect 33197 96389 33243 96435
rect 33321 96389 33367 96435
rect 33445 96389 33491 96435
rect 33569 96389 33615 96435
rect 33693 96389 33739 96435
rect 33817 96389 33863 96435
rect 33941 96389 33987 96435
rect 34065 96389 34111 96435
rect 34189 96389 34235 96435
rect 34313 96389 34359 96435
rect 34437 96389 34483 96435
rect 34561 96389 34607 96435
rect 34685 96389 34731 96435
rect 34809 96389 34855 96435
rect 34933 96389 34979 96435
rect 35057 96389 35103 96435
rect 35181 96389 35227 96435
rect 35305 96389 35351 96435
rect 35429 96389 35475 96435
rect 35553 96389 35599 96435
rect 35677 96389 35723 96435
rect 35801 96389 35847 96435
rect 35925 96389 35971 96435
rect 36049 96389 36095 96435
rect 36173 96389 36219 96435
rect 36297 96389 36343 96435
rect 36421 96389 36467 96435
rect 36545 96389 36591 96435
rect 36669 96389 36715 96435
rect 36793 96389 36839 96435
rect 36917 96389 36963 96435
rect 37041 96389 37087 96435
rect 37165 96389 37211 96435
rect 37289 96389 37335 96435
rect 37413 96389 37459 96435
rect 37537 96389 37583 96435
rect 37661 96389 37707 96435
rect 37785 96389 37831 96435
rect 37909 96389 37955 96435
rect 38033 96389 38079 96435
rect 38157 96389 38203 96435
rect 38281 96389 38327 96435
rect 38405 96389 38451 96435
rect 38529 96389 38575 96435
rect 38653 96389 38699 96435
rect 38777 96389 38823 96435
rect 38901 96389 38947 96435
rect 39025 96389 39071 96435
rect 39149 96389 39195 96435
rect 39273 96389 39319 96435
rect 39397 96389 39443 96435
rect 39521 96389 39567 96435
rect 39645 96389 39691 96435
rect 39769 96389 39815 96435
rect 39893 96389 39939 96435
rect 40017 96389 40063 96435
rect 40141 96389 40187 96435
rect 40265 96389 40311 96435
rect 40389 96389 40435 96435
rect 40513 96389 40559 96435
rect 40637 96389 40683 96435
rect 40761 96389 40807 96435
rect 40885 96389 40931 96435
rect 41009 96389 41055 96435
rect 41133 96389 41179 96435
rect 41257 96389 41303 96435
rect 41381 96389 41427 96435
rect 41505 96389 41551 96435
rect 41629 96389 41675 96435
rect 41753 96389 41799 96435
rect 41877 96389 41923 96435
rect 42001 96389 42047 96435
rect 42125 96389 42171 96435
rect 42249 96389 42295 96435
rect 42373 96389 42419 96435
rect 42497 96389 42543 96435
rect 42621 96389 42667 96435
rect 42745 96389 42791 96435
rect 42869 96389 42915 96435
rect 42993 96389 43039 96435
rect 43117 96389 43163 96435
rect 43241 96389 43287 96435
rect 43365 96389 43411 96435
rect 43489 96389 43535 96435
rect 43613 96389 43659 96435
rect 43737 96389 43783 96435
rect 43861 96389 43907 96435
rect 43985 96389 44031 96435
rect 44109 96389 44155 96435
rect 44233 96389 44279 96435
rect 44357 96389 44403 96435
rect 44481 96389 44527 96435
rect 44605 96389 44651 96435
rect 44729 96389 44775 96435
rect 44853 96389 44899 96435
rect 44977 96389 45023 96435
rect 45101 96389 45147 96435
rect 45225 96389 45271 96435
rect 45349 96389 45395 96435
rect 45473 96389 45519 96435
rect 45597 96389 45643 96435
rect 45721 96389 45767 96435
rect 45845 96389 45891 96435
rect 45969 96389 46015 96435
rect 46093 96389 46139 96435
rect 46217 96389 46263 96435
rect 46341 96389 46387 96435
rect 46465 96389 46511 96435
rect 46589 96389 46635 96435
rect 46713 96389 46759 96435
rect 46837 96389 46883 96435
rect 46961 96389 47007 96435
rect 47085 96389 47131 96435
rect 47209 96389 47255 96435
rect 47333 96389 47379 96435
rect 47457 96389 47503 96435
rect 47581 96389 47627 96435
rect 47705 96389 47751 96435
rect 47829 96389 47875 96435
rect 47953 96389 47999 96435
rect 48077 96389 48123 96435
rect 48201 96389 48247 96435
rect 48325 96389 48371 96435
rect 48449 96389 48495 96435
rect 48573 96389 48619 96435
rect 48697 96389 48743 96435
rect 48821 96389 48867 96435
rect 48945 96389 48991 96435
rect 49069 96389 49115 96435
rect 49193 96389 49239 96435
rect 49317 96389 49363 96435
rect 49441 96389 49487 96435
rect 49565 96389 49611 96435
rect 49689 96389 49735 96435
rect 49813 96389 49859 96435
rect 49937 96389 49983 96435
rect 50061 96389 50107 96435
rect 50185 96389 50231 96435
rect 50309 96389 50355 96435
rect 50433 96389 50479 96435
rect 50557 96389 50603 96435
rect 50681 96389 50727 96435
rect 50805 96389 50851 96435
rect 50929 96389 50975 96435
rect 51053 96389 51099 96435
rect 51177 96389 51223 96435
rect 51301 96389 51347 96435
rect 51425 96389 51471 96435
rect 51549 96389 51595 96435
rect 51673 96389 51719 96435
rect 51797 96389 51843 96435
rect 51921 96389 51967 96435
rect 52045 96389 52091 96435
rect 52169 96389 52215 96435
rect 52293 96389 52339 96435
rect 52417 96389 52463 96435
rect 52541 96389 52587 96435
rect 52665 96389 52711 96435
rect 52789 96389 52835 96435
rect 52913 96389 52959 96435
rect 53037 96389 53083 96435
rect 53161 96389 53207 96435
rect 53285 96389 53331 96435
rect 53409 96389 53455 96435
rect 53533 96389 53579 96435
rect 53657 96389 53703 96435
rect 53781 96389 53827 96435
rect 53905 96389 53951 96435
rect 54029 96389 54075 96435
rect 54153 96389 54199 96435
rect 54277 96389 54323 96435
rect 54401 96389 54447 96435
rect 54525 96389 54571 96435
rect 54649 96389 54695 96435
rect 54773 96389 54819 96435
rect 54897 96389 54943 96435
rect 55021 96389 55067 96435
rect 55145 96389 55191 96435
rect 55269 96389 55315 96435
rect 55393 96389 55439 96435
rect 55517 96389 55563 96435
rect 55641 96389 55687 96435
rect 55765 96389 55811 96435
rect 55889 96389 55935 96435
rect 56013 96389 56059 96435
rect 56137 96389 56183 96435
rect 56261 96389 56307 96435
rect 56385 96389 56431 96435
rect 56509 96389 56555 96435
rect 56633 96389 56679 96435
rect 56757 96389 56803 96435
rect 56881 96389 56927 96435
rect 57005 96389 57051 96435
rect 57129 96389 57175 96435
rect 57253 96389 57299 96435
rect 57377 96389 57423 96435
rect 57501 96389 57547 96435
rect 57625 96389 57671 96435
rect 57749 96389 57795 96435
rect 57873 96389 57919 96435
rect 57997 96389 58043 96435
rect 58121 96389 58167 96435
rect 58245 96389 58291 96435
rect 58369 96389 58415 96435
rect 58493 96389 58539 96435
rect 58617 96389 58663 96435
rect 58741 96389 58787 96435
rect 58865 96389 58911 96435
rect 58989 96389 59035 96435
rect 59113 96389 59159 96435
rect 59237 96389 59283 96435
rect 59361 96389 59407 96435
rect 59485 96389 59531 96435
rect 59609 96389 59655 96435
rect 59733 96389 59779 96435
rect 59857 96389 59903 96435
rect 59981 96389 60027 96435
rect 60105 96389 60151 96435
rect 60229 96389 60275 96435
rect 60353 96389 60399 96435
rect 60477 96389 60523 96435
rect 60601 96389 60647 96435
rect 60725 96389 60771 96435
rect 60849 96389 60895 96435
rect 60973 96389 61019 96435
rect 61097 96389 61143 96435
rect 61221 96389 61267 96435
rect 61345 96389 61391 96435
rect 61469 96389 61515 96435
rect 61593 96389 61639 96435
rect 61717 96389 61763 96435
rect 61841 96389 61887 96435
rect 61965 96389 62011 96435
rect 62089 96389 62135 96435
rect 62213 96389 62259 96435
rect 62337 96389 62383 96435
rect 62461 96389 62507 96435
rect 62585 96389 62631 96435
rect 62709 96389 62755 96435
rect 62833 96389 62879 96435
rect 62957 96389 63003 96435
rect 63081 96389 63127 96435
rect 63205 96389 63251 96435
rect 63329 96389 63375 96435
rect 63453 96389 63499 96435
rect 63577 96389 63623 96435
rect 63701 96389 63747 96435
rect 63825 96389 63871 96435
rect 63949 96389 63995 96435
rect 64073 96389 64119 96435
rect 64197 96389 64243 96435
rect 64321 96389 64367 96435
rect 64445 96389 64491 96435
rect 64569 96389 64615 96435
rect 64693 96389 64739 96435
rect 64817 96389 64863 96435
rect 64941 96389 64987 96435
rect 65065 96389 65111 96435
rect 65189 96389 65235 96435
rect 65313 96389 65359 96435
rect 65437 96389 65483 96435
rect 65561 96389 65607 96435
rect 65685 96389 65731 96435
rect 65809 96389 65855 96435
rect 65933 96389 65979 96435
rect 66057 96389 66103 96435
rect 66181 96389 66227 96435
rect 66305 96389 66351 96435
rect 66429 96389 66475 96435
rect 66553 96389 66599 96435
rect 66677 96389 66723 96435
rect 66801 96389 66847 96435
rect 66925 96389 66971 96435
rect 67049 96389 67095 96435
rect 67173 96389 67219 96435
rect 67297 96389 67343 96435
rect 67421 96389 67467 96435
rect 67545 96389 67591 96435
rect 67669 96389 67715 96435
rect 67793 96389 67839 96435
rect 67917 96389 67963 96435
rect 68041 96389 68087 96435
rect 68165 96389 68211 96435
rect 68289 96389 68335 96435
rect 68413 96389 68459 96435
rect 68537 96389 68583 96435
rect 68661 96389 68707 96435
rect 68785 96389 68831 96435
rect 68909 96389 68955 96435
rect 69033 96389 69079 96435
rect 69157 96389 69203 96435
rect 69281 96389 69327 96435
rect 69405 96389 69451 96435
rect 69529 96389 69575 96435
rect 69653 96389 69699 96435
rect 69777 96389 69823 96435
rect 69901 96389 69947 96435
rect 70025 96389 70071 96435
rect 70149 96389 70195 96435
rect 70273 96389 70319 96435
rect 70397 96389 70443 96435
rect 70521 96389 70567 96435
rect 70645 96389 70691 96435
rect 70769 96389 70815 96435
rect 70893 96389 70939 96435
rect 71017 96389 71063 96435
rect 71141 96389 71187 96435
rect 71265 96389 71311 96435
rect 71389 96389 71435 96435
rect 71513 96389 71559 96435
rect 71637 96389 71683 96435
rect 71761 96389 71807 96435
rect 71885 96389 71931 96435
rect 72009 96389 72055 96435
rect 72133 96389 72179 96435
rect 72257 96389 72303 96435
rect 72381 96389 72427 96435
rect 72505 96389 72551 96435
rect 72629 96389 72675 96435
rect 72753 96389 72799 96435
rect 72877 96389 72923 96435
rect 73001 96389 73047 96435
rect 73125 96389 73171 96435
rect 73249 96389 73295 96435
rect 73373 96389 73419 96435
rect 73497 96389 73543 96435
rect 73621 96389 73667 96435
rect 73745 96389 73791 96435
rect 73869 96389 73915 96435
rect 73993 96389 74039 96435
rect 74117 96389 74163 96435
rect 74241 96389 74287 96435
rect 74365 96389 74411 96435
rect 74489 96389 74535 96435
rect 74613 96389 74659 96435
rect 74737 96389 74783 96435
rect 74861 96389 74907 96435
rect 74985 96389 75031 96435
rect 75109 96389 75155 96435
rect 75233 96389 75279 96435
rect 75357 96389 75403 96435
rect 75481 96389 75527 96435
rect 75605 96389 75651 96435
rect 75729 96389 75775 96435
rect 75853 96389 75899 96435
rect 75977 96389 76023 96435
rect 76101 96389 76147 96435
rect 76225 96389 76271 96435
rect 76349 96389 76395 96435
rect 76473 96389 76519 96435
rect 76597 96389 76643 96435
rect 76721 96389 76767 96435
rect 76845 96389 76891 96435
rect 76969 96389 77015 96435
rect 77093 96389 77139 96435
rect 77217 96389 77263 96435
rect 77341 96389 77387 96435
rect 77465 96389 77511 96435
rect 77589 96389 77635 96435
rect 77713 96389 77759 96435
rect 77837 96389 77883 96435
rect 77961 96389 78007 96435
rect 78085 96389 78131 96435
rect 78209 96389 78255 96435
rect 78333 96389 78379 96435
rect 78457 96389 78503 96435
rect 78581 96389 78627 96435
rect 78705 96389 78751 96435
rect 78829 96389 78875 96435
rect 78953 96389 78999 96435
rect 79077 96389 79123 96435
rect 79201 96389 79247 96435
rect 79325 96389 79371 96435
rect 79449 96389 79495 96435
rect 79573 96389 79619 96435
rect 79697 96389 79743 96435
rect 79821 96389 79867 96435
rect 79945 96389 79991 96435
rect 80069 96389 80115 96435
rect 80193 96389 80239 96435
rect 80317 96389 80363 96435
rect 80441 96389 80487 96435
rect 80565 96389 80611 96435
rect 80689 96389 80735 96435
rect 80813 96389 80859 96435
rect 80937 96389 80983 96435
rect 81061 96389 81107 96435
rect 81185 96389 81231 96435
rect 81309 96389 81355 96435
rect 81433 96389 81479 96435
rect 81557 96389 81603 96435
rect 81681 96389 81727 96435
rect 81805 96389 81851 96435
rect 81929 96389 81975 96435
rect 82053 96389 82099 96435
rect 82177 96389 82223 96435
rect 82301 96389 82347 96435
rect 82425 96389 82471 96435
rect 82549 96389 82595 96435
rect 82673 96389 82719 96435
rect 82797 96389 82843 96435
rect 82921 96389 82967 96435
rect 83045 96389 83091 96435
rect 83169 96389 83215 96435
rect 83293 96389 83339 96435
rect 83417 96389 83463 96435
rect 83541 96389 83587 96435
rect 83665 96389 83711 96435
rect 83789 96389 83835 96435
rect 83913 96389 83959 96435
rect 84037 96389 84083 96435
rect 84161 96389 84207 96435
rect 84285 96389 84331 96435
rect 84409 96389 84455 96435
rect 84533 96389 84579 96435
rect 84657 96389 84703 96435
rect 84781 96389 84827 96435
rect 84905 96389 84951 96435
rect 85029 96389 85075 96435
rect 85153 96389 85199 96435
rect 85277 96389 85323 96435
rect 85401 96389 85447 96435
rect 85525 96389 85571 96435
rect 85649 96389 85695 96435
rect 89 96265 135 96311
rect 213 96265 259 96311
rect 337 96265 383 96311
rect 461 96265 507 96311
rect 585 96265 631 96311
rect 709 96265 755 96311
rect 833 96265 879 96311
rect 957 96265 1003 96311
rect 1081 96265 1127 96311
rect 1205 96265 1251 96311
rect 1329 96265 1375 96311
rect 1453 96265 1499 96311
rect 1577 96265 1623 96311
rect 1701 96265 1747 96311
rect 1825 96265 1871 96311
rect 1949 96265 1995 96311
rect 2073 96265 2119 96311
rect 2197 96265 2243 96311
rect 2321 96265 2367 96311
rect 2445 96265 2491 96311
rect 2569 96265 2615 96311
rect 2693 96265 2739 96311
rect 2817 96265 2863 96311
rect 2941 96265 2987 96311
rect 3065 96265 3111 96311
rect 3189 96265 3235 96311
rect 3313 96265 3359 96311
rect 3437 96265 3483 96311
rect 3561 96265 3607 96311
rect 3685 96265 3731 96311
rect 3809 96265 3855 96311
rect 3933 96265 3979 96311
rect 4057 96265 4103 96311
rect 4181 96265 4227 96311
rect 4305 96265 4351 96311
rect 4429 96265 4475 96311
rect 4553 96265 4599 96311
rect 4677 96265 4723 96311
rect 4801 96265 4847 96311
rect 4925 96265 4971 96311
rect 5049 96265 5095 96311
rect 5173 96265 5219 96311
rect 5297 96265 5343 96311
rect 5421 96265 5467 96311
rect 5545 96265 5591 96311
rect 5669 96265 5715 96311
rect 5793 96265 5839 96311
rect 5917 96265 5963 96311
rect 6041 96265 6087 96311
rect 6165 96265 6211 96311
rect 6289 96265 6335 96311
rect 6413 96265 6459 96311
rect 6537 96265 6583 96311
rect 6661 96265 6707 96311
rect 6785 96265 6831 96311
rect 6909 96265 6955 96311
rect 7033 96265 7079 96311
rect 7157 96265 7203 96311
rect 7281 96265 7327 96311
rect 7405 96265 7451 96311
rect 7529 96265 7575 96311
rect 7653 96265 7699 96311
rect 7777 96265 7823 96311
rect 7901 96265 7947 96311
rect 8025 96265 8071 96311
rect 8149 96265 8195 96311
rect 8273 96265 8319 96311
rect 8397 96265 8443 96311
rect 8521 96265 8567 96311
rect 8645 96265 8691 96311
rect 8769 96265 8815 96311
rect 8893 96265 8939 96311
rect 9017 96265 9063 96311
rect 9141 96265 9187 96311
rect 9265 96265 9311 96311
rect 9389 96265 9435 96311
rect 9513 96265 9559 96311
rect 9637 96265 9683 96311
rect 9761 96265 9807 96311
rect 9885 96265 9931 96311
rect 10009 96265 10055 96311
rect 10133 96265 10179 96311
rect 10257 96265 10303 96311
rect 10381 96265 10427 96311
rect 10505 96265 10551 96311
rect 10629 96265 10675 96311
rect 10753 96265 10799 96311
rect 10877 96265 10923 96311
rect 11001 96265 11047 96311
rect 11125 96265 11171 96311
rect 11249 96265 11295 96311
rect 11373 96265 11419 96311
rect 11497 96265 11543 96311
rect 11621 96265 11667 96311
rect 11745 96265 11791 96311
rect 11869 96265 11915 96311
rect 11993 96265 12039 96311
rect 12117 96265 12163 96311
rect 12241 96265 12287 96311
rect 12365 96265 12411 96311
rect 12489 96265 12535 96311
rect 12613 96265 12659 96311
rect 12737 96265 12783 96311
rect 12861 96265 12907 96311
rect 12985 96265 13031 96311
rect 13109 96265 13155 96311
rect 13233 96265 13279 96311
rect 13357 96265 13403 96311
rect 13481 96265 13527 96311
rect 13605 96265 13651 96311
rect 13729 96265 13775 96311
rect 13853 96265 13899 96311
rect 13977 96265 14023 96311
rect 14101 96265 14147 96311
rect 14225 96265 14271 96311
rect 14349 96265 14395 96311
rect 14473 96265 14519 96311
rect 14597 96265 14643 96311
rect 14721 96265 14767 96311
rect 14845 96265 14891 96311
rect 14969 96265 15015 96311
rect 15093 96265 15139 96311
rect 15217 96265 15263 96311
rect 15341 96265 15387 96311
rect 15465 96265 15511 96311
rect 15589 96265 15635 96311
rect 15713 96265 15759 96311
rect 15837 96265 15883 96311
rect 15961 96265 16007 96311
rect 16085 96265 16131 96311
rect 16209 96265 16255 96311
rect 16333 96265 16379 96311
rect 16457 96265 16503 96311
rect 16581 96265 16627 96311
rect 16705 96265 16751 96311
rect 16829 96265 16875 96311
rect 16953 96265 16999 96311
rect 17077 96265 17123 96311
rect 17201 96265 17247 96311
rect 17325 96265 17371 96311
rect 17449 96265 17495 96311
rect 17573 96265 17619 96311
rect 17697 96265 17743 96311
rect 17821 96265 17867 96311
rect 17945 96265 17991 96311
rect 18069 96265 18115 96311
rect 18193 96265 18239 96311
rect 18317 96265 18363 96311
rect 18441 96265 18487 96311
rect 18565 96265 18611 96311
rect 18689 96265 18735 96311
rect 18813 96265 18859 96311
rect 18937 96265 18983 96311
rect 19061 96265 19107 96311
rect 19185 96265 19231 96311
rect 19309 96265 19355 96311
rect 19433 96265 19479 96311
rect 19557 96265 19603 96311
rect 19681 96265 19727 96311
rect 19805 96265 19851 96311
rect 19929 96265 19975 96311
rect 20053 96265 20099 96311
rect 20177 96265 20223 96311
rect 20301 96265 20347 96311
rect 20425 96265 20471 96311
rect 20549 96265 20595 96311
rect 20673 96265 20719 96311
rect 20797 96265 20843 96311
rect 20921 96265 20967 96311
rect 21045 96265 21091 96311
rect 21169 96265 21215 96311
rect 21293 96265 21339 96311
rect 21417 96265 21463 96311
rect 21541 96265 21587 96311
rect 21665 96265 21711 96311
rect 21789 96265 21835 96311
rect 21913 96265 21959 96311
rect 22037 96265 22083 96311
rect 22161 96265 22207 96311
rect 22285 96265 22331 96311
rect 22409 96265 22455 96311
rect 22533 96265 22579 96311
rect 22657 96265 22703 96311
rect 22781 96265 22827 96311
rect 22905 96265 22951 96311
rect 23029 96265 23075 96311
rect 23153 96265 23199 96311
rect 23277 96265 23323 96311
rect 23401 96265 23447 96311
rect 23525 96265 23571 96311
rect 23649 96265 23695 96311
rect 23773 96265 23819 96311
rect 23897 96265 23943 96311
rect 24021 96265 24067 96311
rect 24145 96265 24191 96311
rect 24269 96265 24315 96311
rect 24393 96265 24439 96311
rect 24517 96265 24563 96311
rect 24641 96265 24687 96311
rect 24765 96265 24811 96311
rect 24889 96265 24935 96311
rect 25013 96265 25059 96311
rect 25137 96265 25183 96311
rect 25261 96265 25307 96311
rect 25385 96265 25431 96311
rect 25509 96265 25555 96311
rect 25633 96265 25679 96311
rect 25757 96265 25803 96311
rect 25881 96265 25927 96311
rect 26005 96265 26051 96311
rect 26129 96265 26175 96311
rect 26253 96265 26299 96311
rect 26377 96265 26423 96311
rect 26501 96265 26547 96311
rect 26625 96265 26671 96311
rect 26749 96265 26795 96311
rect 26873 96265 26919 96311
rect 26997 96265 27043 96311
rect 27121 96265 27167 96311
rect 27245 96265 27291 96311
rect 27369 96265 27415 96311
rect 27493 96265 27539 96311
rect 27617 96265 27663 96311
rect 27741 96265 27787 96311
rect 27865 96265 27911 96311
rect 27989 96265 28035 96311
rect 28113 96265 28159 96311
rect 28237 96265 28283 96311
rect 28361 96265 28407 96311
rect 28485 96265 28531 96311
rect 28609 96265 28655 96311
rect 28733 96265 28779 96311
rect 28857 96265 28903 96311
rect 28981 96265 29027 96311
rect 29105 96265 29151 96311
rect 29229 96265 29275 96311
rect 29353 96265 29399 96311
rect 29477 96265 29523 96311
rect 29601 96265 29647 96311
rect 29725 96265 29771 96311
rect 29849 96265 29895 96311
rect 29973 96265 30019 96311
rect 30097 96265 30143 96311
rect 30221 96265 30267 96311
rect 30345 96265 30391 96311
rect 30469 96265 30515 96311
rect 30593 96265 30639 96311
rect 30717 96265 30763 96311
rect 30841 96265 30887 96311
rect 30965 96265 31011 96311
rect 31089 96265 31135 96311
rect 31213 96265 31259 96311
rect 31337 96265 31383 96311
rect 31461 96265 31507 96311
rect 31585 96265 31631 96311
rect 31709 96265 31755 96311
rect 31833 96265 31879 96311
rect 31957 96265 32003 96311
rect 32081 96265 32127 96311
rect 32205 96265 32251 96311
rect 32329 96265 32375 96311
rect 32453 96265 32499 96311
rect 32577 96265 32623 96311
rect 32701 96265 32747 96311
rect 32825 96265 32871 96311
rect 32949 96265 32995 96311
rect 33073 96265 33119 96311
rect 33197 96265 33243 96311
rect 33321 96265 33367 96311
rect 33445 96265 33491 96311
rect 33569 96265 33615 96311
rect 33693 96265 33739 96311
rect 33817 96265 33863 96311
rect 33941 96265 33987 96311
rect 34065 96265 34111 96311
rect 34189 96265 34235 96311
rect 34313 96265 34359 96311
rect 34437 96265 34483 96311
rect 34561 96265 34607 96311
rect 34685 96265 34731 96311
rect 34809 96265 34855 96311
rect 34933 96265 34979 96311
rect 35057 96265 35103 96311
rect 35181 96265 35227 96311
rect 35305 96265 35351 96311
rect 35429 96265 35475 96311
rect 35553 96265 35599 96311
rect 35677 96265 35723 96311
rect 35801 96265 35847 96311
rect 35925 96265 35971 96311
rect 36049 96265 36095 96311
rect 36173 96265 36219 96311
rect 36297 96265 36343 96311
rect 36421 96265 36467 96311
rect 36545 96265 36591 96311
rect 36669 96265 36715 96311
rect 36793 96265 36839 96311
rect 36917 96265 36963 96311
rect 37041 96265 37087 96311
rect 37165 96265 37211 96311
rect 37289 96265 37335 96311
rect 37413 96265 37459 96311
rect 37537 96265 37583 96311
rect 37661 96265 37707 96311
rect 37785 96265 37831 96311
rect 37909 96265 37955 96311
rect 38033 96265 38079 96311
rect 38157 96265 38203 96311
rect 38281 96265 38327 96311
rect 38405 96265 38451 96311
rect 38529 96265 38575 96311
rect 38653 96265 38699 96311
rect 38777 96265 38823 96311
rect 38901 96265 38947 96311
rect 39025 96265 39071 96311
rect 39149 96265 39195 96311
rect 39273 96265 39319 96311
rect 39397 96265 39443 96311
rect 39521 96265 39567 96311
rect 39645 96265 39691 96311
rect 39769 96265 39815 96311
rect 39893 96265 39939 96311
rect 40017 96265 40063 96311
rect 40141 96265 40187 96311
rect 40265 96265 40311 96311
rect 40389 96265 40435 96311
rect 40513 96265 40559 96311
rect 40637 96265 40683 96311
rect 40761 96265 40807 96311
rect 40885 96265 40931 96311
rect 41009 96265 41055 96311
rect 41133 96265 41179 96311
rect 41257 96265 41303 96311
rect 41381 96265 41427 96311
rect 41505 96265 41551 96311
rect 41629 96265 41675 96311
rect 41753 96265 41799 96311
rect 41877 96265 41923 96311
rect 42001 96265 42047 96311
rect 42125 96265 42171 96311
rect 42249 96265 42295 96311
rect 42373 96265 42419 96311
rect 42497 96265 42543 96311
rect 42621 96265 42667 96311
rect 42745 96265 42791 96311
rect 42869 96265 42915 96311
rect 42993 96265 43039 96311
rect 43117 96265 43163 96311
rect 43241 96265 43287 96311
rect 43365 96265 43411 96311
rect 43489 96265 43535 96311
rect 43613 96265 43659 96311
rect 43737 96265 43783 96311
rect 43861 96265 43907 96311
rect 43985 96265 44031 96311
rect 44109 96265 44155 96311
rect 44233 96265 44279 96311
rect 44357 96265 44403 96311
rect 44481 96265 44527 96311
rect 44605 96265 44651 96311
rect 44729 96265 44775 96311
rect 44853 96265 44899 96311
rect 44977 96265 45023 96311
rect 45101 96265 45147 96311
rect 45225 96265 45271 96311
rect 45349 96265 45395 96311
rect 45473 96265 45519 96311
rect 45597 96265 45643 96311
rect 45721 96265 45767 96311
rect 45845 96265 45891 96311
rect 45969 96265 46015 96311
rect 46093 96265 46139 96311
rect 46217 96265 46263 96311
rect 46341 96265 46387 96311
rect 46465 96265 46511 96311
rect 46589 96265 46635 96311
rect 46713 96265 46759 96311
rect 46837 96265 46883 96311
rect 46961 96265 47007 96311
rect 47085 96265 47131 96311
rect 47209 96265 47255 96311
rect 47333 96265 47379 96311
rect 47457 96265 47503 96311
rect 47581 96265 47627 96311
rect 47705 96265 47751 96311
rect 47829 96265 47875 96311
rect 47953 96265 47999 96311
rect 48077 96265 48123 96311
rect 48201 96265 48247 96311
rect 48325 96265 48371 96311
rect 48449 96265 48495 96311
rect 48573 96265 48619 96311
rect 48697 96265 48743 96311
rect 48821 96265 48867 96311
rect 48945 96265 48991 96311
rect 49069 96265 49115 96311
rect 49193 96265 49239 96311
rect 49317 96265 49363 96311
rect 49441 96265 49487 96311
rect 49565 96265 49611 96311
rect 49689 96265 49735 96311
rect 49813 96265 49859 96311
rect 49937 96265 49983 96311
rect 50061 96265 50107 96311
rect 50185 96265 50231 96311
rect 50309 96265 50355 96311
rect 50433 96265 50479 96311
rect 50557 96265 50603 96311
rect 50681 96265 50727 96311
rect 50805 96265 50851 96311
rect 50929 96265 50975 96311
rect 51053 96265 51099 96311
rect 51177 96265 51223 96311
rect 51301 96265 51347 96311
rect 51425 96265 51471 96311
rect 51549 96265 51595 96311
rect 51673 96265 51719 96311
rect 51797 96265 51843 96311
rect 51921 96265 51967 96311
rect 52045 96265 52091 96311
rect 52169 96265 52215 96311
rect 52293 96265 52339 96311
rect 52417 96265 52463 96311
rect 52541 96265 52587 96311
rect 52665 96265 52711 96311
rect 52789 96265 52835 96311
rect 52913 96265 52959 96311
rect 53037 96265 53083 96311
rect 53161 96265 53207 96311
rect 53285 96265 53331 96311
rect 53409 96265 53455 96311
rect 53533 96265 53579 96311
rect 53657 96265 53703 96311
rect 53781 96265 53827 96311
rect 53905 96265 53951 96311
rect 54029 96265 54075 96311
rect 54153 96265 54199 96311
rect 54277 96265 54323 96311
rect 54401 96265 54447 96311
rect 54525 96265 54571 96311
rect 54649 96265 54695 96311
rect 54773 96265 54819 96311
rect 54897 96265 54943 96311
rect 55021 96265 55067 96311
rect 55145 96265 55191 96311
rect 55269 96265 55315 96311
rect 55393 96265 55439 96311
rect 55517 96265 55563 96311
rect 55641 96265 55687 96311
rect 55765 96265 55811 96311
rect 55889 96265 55935 96311
rect 56013 96265 56059 96311
rect 56137 96265 56183 96311
rect 56261 96265 56307 96311
rect 56385 96265 56431 96311
rect 56509 96265 56555 96311
rect 56633 96265 56679 96311
rect 56757 96265 56803 96311
rect 56881 96265 56927 96311
rect 57005 96265 57051 96311
rect 57129 96265 57175 96311
rect 57253 96265 57299 96311
rect 57377 96265 57423 96311
rect 57501 96265 57547 96311
rect 57625 96265 57671 96311
rect 57749 96265 57795 96311
rect 57873 96265 57919 96311
rect 57997 96265 58043 96311
rect 58121 96265 58167 96311
rect 58245 96265 58291 96311
rect 58369 96265 58415 96311
rect 58493 96265 58539 96311
rect 58617 96265 58663 96311
rect 58741 96265 58787 96311
rect 58865 96265 58911 96311
rect 58989 96265 59035 96311
rect 59113 96265 59159 96311
rect 59237 96265 59283 96311
rect 59361 96265 59407 96311
rect 59485 96265 59531 96311
rect 59609 96265 59655 96311
rect 59733 96265 59779 96311
rect 59857 96265 59903 96311
rect 59981 96265 60027 96311
rect 60105 96265 60151 96311
rect 60229 96265 60275 96311
rect 60353 96265 60399 96311
rect 60477 96265 60523 96311
rect 60601 96265 60647 96311
rect 60725 96265 60771 96311
rect 60849 96265 60895 96311
rect 60973 96265 61019 96311
rect 61097 96265 61143 96311
rect 61221 96265 61267 96311
rect 61345 96265 61391 96311
rect 61469 96265 61515 96311
rect 61593 96265 61639 96311
rect 61717 96265 61763 96311
rect 61841 96265 61887 96311
rect 61965 96265 62011 96311
rect 62089 96265 62135 96311
rect 62213 96265 62259 96311
rect 62337 96265 62383 96311
rect 62461 96265 62507 96311
rect 62585 96265 62631 96311
rect 62709 96265 62755 96311
rect 62833 96265 62879 96311
rect 62957 96265 63003 96311
rect 63081 96265 63127 96311
rect 63205 96265 63251 96311
rect 63329 96265 63375 96311
rect 63453 96265 63499 96311
rect 63577 96265 63623 96311
rect 63701 96265 63747 96311
rect 63825 96265 63871 96311
rect 63949 96265 63995 96311
rect 64073 96265 64119 96311
rect 64197 96265 64243 96311
rect 64321 96265 64367 96311
rect 64445 96265 64491 96311
rect 64569 96265 64615 96311
rect 64693 96265 64739 96311
rect 64817 96265 64863 96311
rect 64941 96265 64987 96311
rect 65065 96265 65111 96311
rect 65189 96265 65235 96311
rect 65313 96265 65359 96311
rect 65437 96265 65483 96311
rect 65561 96265 65607 96311
rect 65685 96265 65731 96311
rect 65809 96265 65855 96311
rect 65933 96265 65979 96311
rect 66057 96265 66103 96311
rect 66181 96265 66227 96311
rect 66305 96265 66351 96311
rect 66429 96265 66475 96311
rect 66553 96265 66599 96311
rect 66677 96265 66723 96311
rect 66801 96265 66847 96311
rect 66925 96265 66971 96311
rect 67049 96265 67095 96311
rect 67173 96265 67219 96311
rect 67297 96265 67343 96311
rect 67421 96265 67467 96311
rect 67545 96265 67591 96311
rect 67669 96265 67715 96311
rect 67793 96265 67839 96311
rect 67917 96265 67963 96311
rect 68041 96265 68087 96311
rect 68165 96265 68211 96311
rect 68289 96265 68335 96311
rect 68413 96265 68459 96311
rect 68537 96265 68583 96311
rect 68661 96265 68707 96311
rect 68785 96265 68831 96311
rect 68909 96265 68955 96311
rect 69033 96265 69079 96311
rect 69157 96265 69203 96311
rect 69281 96265 69327 96311
rect 69405 96265 69451 96311
rect 69529 96265 69575 96311
rect 69653 96265 69699 96311
rect 69777 96265 69823 96311
rect 69901 96265 69947 96311
rect 70025 96265 70071 96311
rect 70149 96265 70195 96311
rect 70273 96265 70319 96311
rect 70397 96265 70443 96311
rect 70521 96265 70567 96311
rect 70645 96265 70691 96311
rect 70769 96265 70815 96311
rect 70893 96265 70939 96311
rect 71017 96265 71063 96311
rect 71141 96265 71187 96311
rect 71265 96265 71311 96311
rect 71389 96265 71435 96311
rect 71513 96265 71559 96311
rect 71637 96265 71683 96311
rect 71761 96265 71807 96311
rect 71885 96265 71931 96311
rect 72009 96265 72055 96311
rect 72133 96265 72179 96311
rect 72257 96265 72303 96311
rect 72381 96265 72427 96311
rect 72505 96265 72551 96311
rect 72629 96265 72675 96311
rect 72753 96265 72799 96311
rect 72877 96265 72923 96311
rect 73001 96265 73047 96311
rect 73125 96265 73171 96311
rect 73249 96265 73295 96311
rect 73373 96265 73419 96311
rect 73497 96265 73543 96311
rect 73621 96265 73667 96311
rect 73745 96265 73791 96311
rect 73869 96265 73915 96311
rect 73993 96265 74039 96311
rect 74117 96265 74163 96311
rect 74241 96265 74287 96311
rect 74365 96265 74411 96311
rect 74489 96265 74535 96311
rect 74613 96265 74659 96311
rect 74737 96265 74783 96311
rect 74861 96265 74907 96311
rect 74985 96265 75031 96311
rect 75109 96265 75155 96311
rect 75233 96265 75279 96311
rect 75357 96265 75403 96311
rect 75481 96265 75527 96311
rect 75605 96265 75651 96311
rect 75729 96265 75775 96311
rect 75853 96265 75899 96311
rect 75977 96265 76023 96311
rect 76101 96265 76147 96311
rect 76225 96265 76271 96311
rect 76349 96265 76395 96311
rect 76473 96265 76519 96311
rect 76597 96265 76643 96311
rect 76721 96265 76767 96311
rect 76845 96265 76891 96311
rect 76969 96265 77015 96311
rect 77093 96265 77139 96311
rect 77217 96265 77263 96311
rect 77341 96265 77387 96311
rect 77465 96265 77511 96311
rect 77589 96265 77635 96311
rect 77713 96265 77759 96311
rect 77837 96265 77883 96311
rect 77961 96265 78007 96311
rect 78085 96265 78131 96311
rect 78209 96265 78255 96311
rect 78333 96265 78379 96311
rect 78457 96265 78503 96311
rect 78581 96265 78627 96311
rect 78705 96265 78751 96311
rect 78829 96265 78875 96311
rect 78953 96265 78999 96311
rect 79077 96265 79123 96311
rect 79201 96265 79247 96311
rect 79325 96265 79371 96311
rect 79449 96265 79495 96311
rect 79573 96265 79619 96311
rect 79697 96265 79743 96311
rect 79821 96265 79867 96311
rect 79945 96265 79991 96311
rect 80069 96265 80115 96311
rect 80193 96265 80239 96311
rect 80317 96265 80363 96311
rect 80441 96265 80487 96311
rect 80565 96265 80611 96311
rect 80689 96265 80735 96311
rect 80813 96265 80859 96311
rect 80937 96265 80983 96311
rect 81061 96265 81107 96311
rect 81185 96265 81231 96311
rect 81309 96265 81355 96311
rect 81433 96265 81479 96311
rect 81557 96265 81603 96311
rect 81681 96265 81727 96311
rect 81805 96265 81851 96311
rect 81929 96265 81975 96311
rect 82053 96265 82099 96311
rect 82177 96265 82223 96311
rect 82301 96265 82347 96311
rect 82425 96265 82471 96311
rect 82549 96265 82595 96311
rect 82673 96265 82719 96311
rect 82797 96265 82843 96311
rect 82921 96265 82967 96311
rect 83045 96265 83091 96311
rect 83169 96265 83215 96311
rect 83293 96265 83339 96311
rect 83417 96265 83463 96311
rect 83541 96265 83587 96311
rect 83665 96265 83711 96311
rect 83789 96265 83835 96311
rect 83913 96265 83959 96311
rect 84037 96265 84083 96311
rect 84161 96265 84207 96311
rect 84285 96265 84331 96311
rect 84409 96265 84455 96311
rect 84533 96265 84579 96311
rect 84657 96265 84703 96311
rect 84781 96265 84827 96311
rect 84905 96265 84951 96311
rect 85029 96265 85075 96311
rect 85153 96265 85199 96311
rect 85277 96265 85323 96311
rect 85401 96265 85447 96311
rect 85525 96265 85571 96311
rect 85649 96265 85695 96311
rect 89 1117 435 96163
rect 27116 1117 27462 96163
rect 27540 35996 28386 96142
rect 56100 35996 56946 96142
rect 27540 34174 56886 34620
rect 57024 1117 57370 96163
rect 85451 1117 85797 96163
rect 89 969 135 1015
rect 213 969 259 1015
rect 337 969 383 1015
rect 461 969 507 1015
rect 585 969 631 1015
rect 709 969 755 1015
rect 833 969 879 1015
rect 957 969 1003 1015
rect 1081 969 1127 1015
rect 1205 969 1251 1015
rect 1329 969 1375 1015
rect 1453 969 1499 1015
rect 1577 969 1623 1015
rect 1701 969 1747 1015
rect 1825 969 1871 1015
rect 1949 969 1995 1015
rect 2073 969 2119 1015
rect 2197 969 2243 1015
rect 2321 969 2367 1015
rect 2445 969 2491 1015
rect 2569 969 2615 1015
rect 2693 969 2739 1015
rect 2817 969 2863 1015
rect 2941 969 2987 1015
rect 3065 969 3111 1015
rect 3189 969 3235 1015
rect 3313 969 3359 1015
rect 3437 969 3483 1015
rect 3561 969 3607 1015
rect 3685 969 3731 1015
rect 3809 969 3855 1015
rect 3933 969 3979 1015
rect 4057 969 4103 1015
rect 4181 969 4227 1015
rect 4305 969 4351 1015
rect 4429 969 4475 1015
rect 4553 969 4599 1015
rect 4677 969 4723 1015
rect 4801 969 4847 1015
rect 4925 969 4971 1015
rect 5049 969 5095 1015
rect 5173 969 5219 1015
rect 5297 969 5343 1015
rect 5421 969 5467 1015
rect 5545 969 5591 1015
rect 5669 969 5715 1015
rect 5793 969 5839 1015
rect 5917 969 5963 1015
rect 6041 969 6087 1015
rect 6165 969 6211 1015
rect 6289 969 6335 1015
rect 6413 969 6459 1015
rect 6537 969 6583 1015
rect 6661 969 6707 1015
rect 6785 969 6831 1015
rect 6909 969 6955 1015
rect 7033 969 7079 1015
rect 7157 969 7203 1015
rect 7281 969 7327 1015
rect 7405 969 7451 1015
rect 7529 969 7575 1015
rect 7653 969 7699 1015
rect 7777 969 7823 1015
rect 7901 969 7947 1015
rect 8025 969 8071 1015
rect 8149 969 8195 1015
rect 8273 969 8319 1015
rect 8397 969 8443 1015
rect 8521 969 8567 1015
rect 8645 969 8691 1015
rect 8769 969 8815 1015
rect 8893 969 8939 1015
rect 9017 969 9063 1015
rect 9141 969 9187 1015
rect 9265 969 9311 1015
rect 9389 969 9435 1015
rect 9513 969 9559 1015
rect 9637 969 9683 1015
rect 9761 969 9807 1015
rect 9885 969 9931 1015
rect 10009 969 10055 1015
rect 10133 969 10179 1015
rect 10257 969 10303 1015
rect 10381 969 10427 1015
rect 10505 969 10551 1015
rect 10629 969 10675 1015
rect 10753 969 10799 1015
rect 10877 969 10923 1015
rect 11001 969 11047 1015
rect 11125 969 11171 1015
rect 11249 969 11295 1015
rect 11373 969 11419 1015
rect 11497 969 11543 1015
rect 11621 969 11667 1015
rect 11745 969 11791 1015
rect 11869 969 11915 1015
rect 11993 969 12039 1015
rect 12117 969 12163 1015
rect 12241 969 12287 1015
rect 12365 969 12411 1015
rect 12489 969 12535 1015
rect 12613 969 12659 1015
rect 12737 969 12783 1015
rect 12861 969 12907 1015
rect 12985 969 13031 1015
rect 13109 969 13155 1015
rect 13233 969 13279 1015
rect 13357 969 13403 1015
rect 13481 969 13527 1015
rect 13605 969 13651 1015
rect 13729 969 13775 1015
rect 13853 969 13899 1015
rect 13977 969 14023 1015
rect 14101 969 14147 1015
rect 14225 969 14271 1015
rect 14349 969 14395 1015
rect 14473 969 14519 1015
rect 14597 969 14643 1015
rect 14721 969 14767 1015
rect 14845 969 14891 1015
rect 14969 969 15015 1015
rect 15093 969 15139 1015
rect 15217 969 15263 1015
rect 15341 969 15387 1015
rect 15465 969 15511 1015
rect 15589 969 15635 1015
rect 15713 969 15759 1015
rect 15837 969 15883 1015
rect 15961 969 16007 1015
rect 16085 969 16131 1015
rect 16209 969 16255 1015
rect 16333 969 16379 1015
rect 16457 969 16503 1015
rect 16581 969 16627 1015
rect 16705 969 16751 1015
rect 16829 969 16875 1015
rect 16953 969 16999 1015
rect 17077 969 17123 1015
rect 17201 969 17247 1015
rect 17325 969 17371 1015
rect 17449 969 17495 1015
rect 17573 969 17619 1015
rect 17697 969 17743 1015
rect 17821 969 17867 1015
rect 17945 969 17991 1015
rect 18069 969 18115 1015
rect 18193 969 18239 1015
rect 18317 969 18363 1015
rect 18441 969 18487 1015
rect 18565 969 18611 1015
rect 18689 969 18735 1015
rect 18813 969 18859 1015
rect 18937 969 18983 1015
rect 19061 969 19107 1015
rect 19185 969 19231 1015
rect 19309 969 19355 1015
rect 19433 969 19479 1015
rect 19557 969 19603 1015
rect 19681 969 19727 1015
rect 19805 969 19851 1015
rect 19929 969 19975 1015
rect 20053 969 20099 1015
rect 20177 969 20223 1015
rect 20301 969 20347 1015
rect 20425 969 20471 1015
rect 20549 969 20595 1015
rect 20673 969 20719 1015
rect 20797 969 20843 1015
rect 20921 969 20967 1015
rect 21045 969 21091 1015
rect 21169 969 21215 1015
rect 21293 969 21339 1015
rect 21417 969 21463 1015
rect 21541 969 21587 1015
rect 21665 969 21711 1015
rect 21789 969 21835 1015
rect 21913 969 21959 1015
rect 22037 969 22083 1015
rect 22161 969 22207 1015
rect 22285 969 22331 1015
rect 22409 969 22455 1015
rect 22533 969 22579 1015
rect 22657 969 22703 1015
rect 22781 969 22827 1015
rect 22905 969 22951 1015
rect 23029 969 23075 1015
rect 23153 969 23199 1015
rect 23277 969 23323 1015
rect 23401 969 23447 1015
rect 23525 969 23571 1015
rect 23649 969 23695 1015
rect 23773 969 23819 1015
rect 23897 969 23943 1015
rect 24021 969 24067 1015
rect 24145 969 24191 1015
rect 24269 969 24315 1015
rect 24393 969 24439 1015
rect 24517 969 24563 1015
rect 24641 969 24687 1015
rect 24765 969 24811 1015
rect 24889 969 24935 1015
rect 25013 969 25059 1015
rect 25137 969 25183 1015
rect 25261 969 25307 1015
rect 25385 969 25431 1015
rect 25509 969 25555 1015
rect 25633 969 25679 1015
rect 25757 969 25803 1015
rect 25881 969 25927 1015
rect 26005 969 26051 1015
rect 26129 969 26175 1015
rect 26253 969 26299 1015
rect 26377 969 26423 1015
rect 26501 969 26547 1015
rect 26625 969 26671 1015
rect 26749 969 26795 1015
rect 26873 969 26919 1015
rect 26997 969 27043 1015
rect 27121 969 27167 1015
rect 27245 969 27291 1015
rect 27369 969 27415 1015
rect 27493 969 27539 1015
rect 27617 969 27663 1015
rect 27741 969 27787 1015
rect 27865 969 27911 1015
rect 27989 969 28035 1015
rect 28113 969 28159 1015
rect 28237 969 28283 1015
rect 28361 969 28407 1015
rect 28485 969 28531 1015
rect 28609 969 28655 1015
rect 28733 969 28779 1015
rect 28857 969 28903 1015
rect 28981 969 29027 1015
rect 29105 969 29151 1015
rect 29229 969 29275 1015
rect 29353 969 29399 1015
rect 29477 969 29523 1015
rect 29601 969 29647 1015
rect 29725 969 29771 1015
rect 29849 969 29895 1015
rect 29973 969 30019 1015
rect 30097 969 30143 1015
rect 30221 969 30267 1015
rect 30345 969 30391 1015
rect 30469 969 30515 1015
rect 30593 969 30639 1015
rect 30717 969 30763 1015
rect 30841 969 30887 1015
rect 30965 969 31011 1015
rect 31089 969 31135 1015
rect 31213 969 31259 1015
rect 31337 969 31383 1015
rect 31461 969 31507 1015
rect 31585 969 31631 1015
rect 31709 969 31755 1015
rect 31833 969 31879 1015
rect 31957 969 32003 1015
rect 32081 969 32127 1015
rect 32205 969 32251 1015
rect 32329 969 32375 1015
rect 32453 969 32499 1015
rect 32577 969 32623 1015
rect 32701 969 32747 1015
rect 32825 969 32871 1015
rect 32949 969 32995 1015
rect 33073 969 33119 1015
rect 33197 969 33243 1015
rect 33321 969 33367 1015
rect 33445 969 33491 1015
rect 33569 969 33615 1015
rect 33693 969 33739 1015
rect 33817 969 33863 1015
rect 33941 969 33987 1015
rect 34065 969 34111 1015
rect 34189 969 34235 1015
rect 34313 969 34359 1015
rect 34437 969 34483 1015
rect 34561 969 34607 1015
rect 34685 969 34731 1015
rect 34809 969 34855 1015
rect 34933 969 34979 1015
rect 35057 969 35103 1015
rect 35181 969 35227 1015
rect 35305 969 35351 1015
rect 35429 969 35475 1015
rect 35553 969 35599 1015
rect 35677 969 35723 1015
rect 35801 969 35847 1015
rect 35925 969 35971 1015
rect 36049 969 36095 1015
rect 36173 969 36219 1015
rect 36297 969 36343 1015
rect 36421 969 36467 1015
rect 36545 969 36591 1015
rect 36669 969 36715 1015
rect 36793 969 36839 1015
rect 36917 969 36963 1015
rect 37041 969 37087 1015
rect 37165 969 37211 1015
rect 37289 969 37335 1015
rect 37413 969 37459 1015
rect 37537 969 37583 1015
rect 37661 969 37707 1015
rect 37785 969 37831 1015
rect 37909 969 37955 1015
rect 38033 969 38079 1015
rect 38157 969 38203 1015
rect 38281 969 38327 1015
rect 38405 969 38451 1015
rect 38529 969 38575 1015
rect 38653 969 38699 1015
rect 38777 969 38823 1015
rect 38901 969 38947 1015
rect 39025 969 39071 1015
rect 39149 969 39195 1015
rect 39273 969 39319 1015
rect 39397 969 39443 1015
rect 39521 969 39567 1015
rect 39645 969 39691 1015
rect 39769 969 39815 1015
rect 39893 969 39939 1015
rect 40017 969 40063 1015
rect 40141 969 40187 1015
rect 40265 969 40311 1015
rect 40389 969 40435 1015
rect 40513 969 40559 1015
rect 40637 969 40683 1015
rect 40761 969 40807 1015
rect 40885 969 40931 1015
rect 41009 969 41055 1015
rect 41133 969 41179 1015
rect 41257 969 41303 1015
rect 41381 969 41427 1015
rect 41505 969 41551 1015
rect 41629 969 41675 1015
rect 41753 969 41799 1015
rect 41877 969 41923 1015
rect 42001 969 42047 1015
rect 42125 969 42171 1015
rect 42249 969 42295 1015
rect 42373 969 42419 1015
rect 42497 969 42543 1015
rect 42621 969 42667 1015
rect 42745 969 42791 1015
rect 42869 969 42915 1015
rect 42993 969 43039 1015
rect 43117 969 43163 1015
rect 43241 969 43287 1015
rect 43365 969 43411 1015
rect 43489 969 43535 1015
rect 43613 969 43659 1015
rect 43737 969 43783 1015
rect 43861 969 43907 1015
rect 43985 969 44031 1015
rect 44109 969 44155 1015
rect 44233 969 44279 1015
rect 44357 969 44403 1015
rect 44481 969 44527 1015
rect 44605 969 44651 1015
rect 44729 969 44775 1015
rect 44853 969 44899 1015
rect 44977 969 45023 1015
rect 45101 969 45147 1015
rect 45225 969 45271 1015
rect 45349 969 45395 1015
rect 45473 969 45519 1015
rect 45597 969 45643 1015
rect 45721 969 45767 1015
rect 45845 969 45891 1015
rect 45969 969 46015 1015
rect 46093 969 46139 1015
rect 46217 969 46263 1015
rect 46341 969 46387 1015
rect 46465 969 46511 1015
rect 46589 969 46635 1015
rect 46713 969 46759 1015
rect 46837 969 46883 1015
rect 46961 969 47007 1015
rect 47085 969 47131 1015
rect 47209 969 47255 1015
rect 47333 969 47379 1015
rect 47457 969 47503 1015
rect 47581 969 47627 1015
rect 47705 969 47751 1015
rect 47829 969 47875 1015
rect 47953 969 47999 1015
rect 48077 969 48123 1015
rect 48201 969 48247 1015
rect 48325 969 48371 1015
rect 48449 969 48495 1015
rect 48573 969 48619 1015
rect 48697 969 48743 1015
rect 48821 969 48867 1015
rect 48945 969 48991 1015
rect 49069 969 49115 1015
rect 49193 969 49239 1015
rect 49317 969 49363 1015
rect 49441 969 49487 1015
rect 49565 969 49611 1015
rect 49689 969 49735 1015
rect 49813 969 49859 1015
rect 49937 969 49983 1015
rect 50061 969 50107 1015
rect 50185 969 50231 1015
rect 50309 969 50355 1015
rect 50433 969 50479 1015
rect 50557 969 50603 1015
rect 50681 969 50727 1015
rect 50805 969 50851 1015
rect 50929 969 50975 1015
rect 51053 969 51099 1015
rect 51177 969 51223 1015
rect 51301 969 51347 1015
rect 51425 969 51471 1015
rect 51549 969 51595 1015
rect 51673 969 51719 1015
rect 51797 969 51843 1015
rect 51921 969 51967 1015
rect 52045 969 52091 1015
rect 52169 969 52215 1015
rect 52293 969 52339 1015
rect 52417 969 52463 1015
rect 52541 969 52587 1015
rect 52665 969 52711 1015
rect 52789 969 52835 1015
rect 52913 969 52959 1015
rect 53037 969 53083 1015
rect 53161 969 53207 1015
rect 53285 969 53331 1015
rect 53409 969 53455 1015
rect 53533 969 53579 1015
rect 53657 969 53703 1015
rect 53781 969 53827 1015
rect 53905 969 53951 1015
rect 54029 969 54075 1015
rect 54153 969 54199 1015
rect 54277 969 54323 1015
rect 54401 969 54447 1015
rect 54525 969 54571 1015
rect 54649 969 54695 1015
rect 54773 969 54819 1015
rect 54897 969 54943 1015
rect 55021 969 55067 1015
rect 55145 969 55191 1015
rect 55269 969 55315 1015
rect 55393 969 55439 1015
rect 55517 969 55563 1015
rect 55641 969 55687 1015
rect 55765 969 55811 1015
rect 55889 969 55935 1015
rect 56013 969 56059 1015
rect 56137 969 56183 1015
rect 56261 969 56307 1015
rect 56385 969 56431 1015
rect 56509 969 56555 1015
rect 56633 969 56679 1015
rect 56757 969 56803 1015
rect 56881 969 56927 1015
rect 57005 969 57051 1015
rect 57129 969 57175 1015
rect 57253 969 57299 1015
rect 57377 969 57423 1015
rect 57501 969 57547 1015
rect 57625 969 57671 1015
rect 57749 969 57795 1015
rect 57873 969 57919 1015
rect 57997 969 58043 1015
rect 58121 969 58167 1015
rect 58245 969 58291 1015
rect 58369 969 58415 1015
rect 58493 969 58539 1015
rect 58617 969 58663 1015
rect 58741 969 58787 1015
rect 58865 969 58911 1015
rect 58989 969 59035 1015
rect 59113 969 59159 1015
rect 59237 969 59283 1015
rect 59361 969 59407 1015
rect 59485 969 59531 1015
rect 59609 969 59655 1015
rect 59733 969 59779 1015
rect 59857 969 59903 1015
rect 59981 969 60027 1015
rect 60105 969 60151 1015
rect 60229 969 60275 1015
rect 60353 969 60399 1015
rect 60477 969 60523 1015
rect 60601 969 60647 1015
rect 60725 969 60771 1015
rect 60849 969 60895 1015
rect 60973 969 61019 1015
rect 61097 969 61143 1015
rect 61221 969 61267 1015
rect 61345 969 61391 1015
rect 61469 969 61515 1015
rect 61593 969 61639 1015
rect 61717 969 61763 1015
rect 61841 969 61887 1015
rect 61965 969 62011 1015
rect 62089 969 62135 1015
rect 62213 969 62259 1015
rect 62337 969 62383 1015
rect 62461 969 62507 1015
rect 62585 969 62631 1015
rect 62709 969 62755 1015
rect 62833 969 62879 1015
rect 62957 969 63003 1015
rect 63081 969 63127 1015
rect 63205 969 63251 1015
rect 63329 969 63375 1015
rect 63453 969 63499 1015
rect 63577 969 63623 1015
rect 63701 969 63747 1015
rect 63825 969 63871 1015
rect 63949 969 63995 1015
rect 64073 969 64119 1015
rect 64197 969 64243 1015
rect 64321 969 64367 1015
rect 64445 969 64491 1015
rect 64569 969 64615 1015
rect 64693 969 64739 1015
rect 64817 969 64863 1015
rect 64941 969 64987 1015
rect 65065 969 65111 1015
rect 65189 969 65235 1015
rect 65313 969 65359 1015
rect 65437 969 65483 1015
rect 65561 969 65607 1015
rect 65685 969 65731 1015
rect 65809 969 65855 1015
rect 65933 969 65979 1015
rect 66057 969 66103 1015
rect 66181 969 66227 1015
rect 66305 969 66351 1015
rect 66429 969 66475 1015
rect 66553 969 66599 1015
rect 66677 969 66723 1015
rect 66801 969 66847 1015
rect 66925 969 66971 1015
rect 67049 969 67095 1015
rect 67173 969 67219 1015
rect 67297 969 67343 1015
rect 67421 969 67467 1015
rect 67545 969 67591 1015
rect 67669 969 67715 1015
rect 67793 969 67839 1015
rect 67917 969 67963 1015
rect 68041 969 68087 1015
rect 68165 969 68211 1015
rect 68289 969 68335 1015
rect 68413 969 68459 1015
rect 68537 969 68583 1015
rect 68661 969 68707 1015
rect 68785 969 68831 1015
rect 68909 969 68955 1015
rect 69033 969 69079 1015
rect 69157 969 69203 1015
rect 69281 969 69327 1015
rect 69405 969 69451 1015
rect 69529 969 69575 1015
rect 69653 969 69699 1015
rect 69777 969 69823 1015
rect 69901 969 69947 1015
rect 70025 969 70071 1015
rect 70149 969 70195 1015
rect 70273 969 70319 1015
rect 70397 969 70443 1015
rect 70521 969 70567 1015
rect 70645 969 70691 1015
rect 70769 969 70815 1015
rect 70893 969 70939 1015
rect 71017 969 71063 1015
rect 71141 969 71187 1015
rect 71265 969 71311 1015
rect 71389 969 71435 1015
rect 71513 969 71559 1015
rect 71637 969 71683 1015
rect 71761 969 71807 1015
rect 71885 969 71931 1015
rect 72009 969 72055 1015
rect 72133 969 72179 1015
rect 72257 969 72303 1015
rect 72381 969 72427 1015
rect 72505 969 72551 1015
rect 72629 969 72675 1015
rect 72753 969 72799 1015
rect 72877 969 72923 1015
rect 73001 969 73047 1015
rect 73125 969 73171 1015
rect 73249 969 73295 1015
rect 73373 969 73419 1015
rect 73497 969 73543 1015
rect 73621 969 73667 1015
rect 73745 969 73791 1015
rect 73869 969 73915 1015
rect 73993 969 74039 1015
rect 74117 969 74163 1015
rect 74241 969 74287 1015
rect 74365 969 74411 1015
rect 74489 969 74535 1015
rect 74613 969 74659 1015
rect 74737 969 74783 1015
rect 74861 969 74907 1015
rect 74985 969 75031 1015
rect 75109 969 75155 1015
rect 75233 969 75279 1015
rect 75357 969 75403 1015
rect 75481 969 75527 1015
rect 75605 969 75651 1015
rect 75729 969 75775 1015
rect 75853 969 75899 1015
rect 75977 969 76023 1015
rect 76101 969 76147 1015
rect 76225 969 76271 1015
rect 76349 969 76395 1015
rect 76473 969 76519 1015
rect 76597 969 76643 1015
rect 76721 969 76767 1015
rect 76845 969 76891 1015
rect 76969 969 77015 1015
rect 77093 969 77139 1015
rect 77217 969 77263 1015
rect 77341 969 77387 1015
rect 77465 969 77511 1015
rect 77589 969 77635 1015
rect 77713 969 77759 1015
rect 77837 969 77883 1015
rect 77961 969 78007 1015
rect 78085 969 78131 1015
rect 78209 969 78255 1015
rect 78333 969 78379 1015
rect 78457 969 78503 1015
rect 78581 969 78627 1015
rect 78705 969 78751 1015
rect 78829 969 78875 1015
rect 78953 969 78999 1015
rect 79077 969 79123 1015
rect 79201 969 79247 1015
rect 79325 969 79371 1015
rect 79449 969 79495 1015
rect 79573 969 79619 1015
rect 79697 969 79743 1015
rect 79821 969 79867 1015
rect 79945 969 79991 1015
rect 80069 969 80115 1015
rect 80193 969 80239 1015
rect 80317 969 80363 1015
rect 80441 969 80487 1015
rect 80565 969 80611 1015
rect 80689 969 80735 1015
rect 80813 969 80859 1015
rect 80937 969 80983 1015
rect 81061 969 81107 1015
rect 81185 969 81231 1015
rect 81309 969 81355 1015
rect 81433 969 81479 1015
rect 81557 969 81603 1015
rect 81681 969 81727 1015
rect 81805 969 81851 1015
rect 81929 969 81975 1015
rect 82053 969 82099 1015
rect 82177 969 82223 1015
rect 82301 969 82347 1015
rect 82425 969 82471 1015
rect 82549 969 82595 1015
rect 82673 969 82719 1015
rect 82797 969 82843 1015
rect 82921 969 82967 1015
rect 83045 969 83091 1015
rect 83169 969 83215 1015
rect 83293 969 83339 1015
rect 83417 969 83463 1015
rect 83541 969 83587 1015
rect 83665 969 83711 1015
rect 83789 969 83835 1015
rect 83913 969 83959 1015
rect 84037 969 84083 1015
rect 84161 969 84207 1015
rect 84285 969 84331 1015
rect 84409 969 84455 1015
rect 84533 969 84579 1015
rect 84657 969 84703 1015
rect 84781 969 84827 1015
rect 84905 969 84951 1015
rect 85029 969 85075 1015
rect 85153 969 85199 1015
rect 85277 969 85323 1015
rect 85401 969 85447 1015
rect 85525 969 85571 1015
rect 85649 969 85695 1015
rect 89 845 135 891
rect 213 845 259 891
rect 337 845 383 891
rect 461 845 507 891
rect 585 845 631 891
rect 709 845 755 891
rect 833 845 879 891
rect 957 845 1003 891
rect 1081 845 1127 891
rect 1205 845 1251 891
rect 1329 845 1375 891
rect 1453 845 1499 891
rect 1577 845 1623 891
rect 1701 845 1747 891
rect 1825 845 1871 891
rect 1949 845 1995 891
rect 2073 845 2119 891
rect 2197 845 2243 891
rect 2321 845 2367 891
rect 2445 845 2491 891
rect 2569 845 2615 891
rect 2693 845 2739 891
rect 2817 845 2863 891
rect 2941 845 2987 891
rect 3065 845 3111 891
rect 3189 845 3235 891
rect 3313 845 3359 891
rect 3437 845 3483 891
rect 3561 845 3607 891
rect 3685 845 3731 891
rect 3809 845 3855 891
rect 3933 845 3979 891
rect 4057 845 4103 891
rect 4181 845 4227 891
rect 4305 845 4351 891
rect 4429 845 4475 891
rect 4553 845 4599 891
rect 4677 845 4723 891
rect 4801 845 4847 891
rect 4925 845 4971 891
rect 5049 845 5095 891
rect 5173 845 5219 891
rect 5297 845 5343 891
rect 5421 845 5467 891
rect 5545 845 5591 891
rect 5669 845 5715 891
rect 5793 845 5839 891
rect 5917 845 5963 891
rect 6041 845 6087 891
rect 6165 845 6211 891
rect 6289 845 6335 891
rect 6413 845 6459 891
rect 6537 845 6583 891
rect 6661 845 6707 891
rect 6785 845 6831 891
rect 6909 845 6955 891
rect 7033 845 7079 891
rect 7157 845 7203 891
rect 7281 845 7327 891
rect 7405 845 7451 891
rect 7529 845 7575 891
rect 7653 845 7699 891
rect 7777 845 7823 891
rect 7901 845 7947 891
rect 8025 845 8071 891
rect 8149 845 8195 891
rect 8273 845 8319 891
rect 8397 845 8443 891
rect 8521 845 8567 891
rect 8645 845 8691 891
rect 8769 845 8815 891
rect 8893 845 8939 891
rect 9017 845 9063 891
rect 9141 845 9187 891
rect 9265 845 9311 891
rect 9389 845 9435 891
rect 9513 845 9559 891
rect 9637 845 9683 891
rect 9761 845 9807 891
rect 9885 845 9931 891
rect 10009 845 10055 891
rect 10133 845 10179 891
rect 10257 845 10303 891
rect 10381 845 10427 891
rect 10505 845 10551 891
rect 10629 845 10675 891
rect 10753 845 10799 891
rect 10877 845 10923 891
rect 11001 845 11047 891
rect 11125 845 11171 891
rect 11249 845 11295 891
rect 11373 845 11419 891
rect 11497 845 11543 891
rect 11621 845 11667 891
rect 11745 845 11791 891
rect 11869 845 11915 891
rect 11993 845 12039 891
rect 12117 845 12163 891
rect 12241 845 12287 891
rect 12365 845 12411 891
rect 12489 845 12535 891
rect 12613 845 12659 891
rect 12737 845 12783 891
rect 12861 845 12907 891
rect 12985 845 13031 891
rect 13109 845 13155 891
rect 13233 845 13279 891
rect 13357 845 13403 891
rect 13481 845 13527 891
rect 13605 845 13651 891
rect 13729 845 13775 891
rect 13853 845 13899 891
rect 13977 845 14023 891
rect 14101 845 14147 891
rect 14225 845 14271 891
rect 14349 845 14395 891
rect 14473 845 14519 891
rect 14597 845 14643 891
rect 14721 845 14767 891
rect 14845 845 14891 891
rect 14969 845 15015 891
rect 15093 845 15139 891
rect 15217 845 15263 891
rect 15341 845 15387 891
rect 15465 845 15511 891
rect 15589 845 15635 891
rect 15713 845 15759 891
rect 15837 845 15883 891
rect 15961 845 16007 891
rect 16085 845 16131 891
rect 16209 845 16255 891
rect 16333 845 16379 891
rect 16457 845 16503 891
rect 16581 845 16627 891
rect 16705 845 16751 891
rect 16829 845 16875 891
rect 16953 845 16999 891
rect 17077 845 17123 891
rect 17201 845 17247 891
rect 17325 845 17371 891
rect 17449 845 17495 891
rect 17573 845 17619 891
rect 17697 845 17743 891
rect 17821 845 17867 891
rect 17945 845 17991 891
rect 18069 845 18115 891
rect 18193 845 18239 891
rect 18317 845 18363 891
rect 18441 845 18487 891
rect 18565 845 18611 891
rect 18689 845 18735 891
rect 18813 845 18859 891
rect 18937 845 18983 891
rect 19061 845 19107 891
rect 19185 845 19231 891
rect 19309 845 19355 891
rect 19433 845 19479 891
rect 19557 845 19603 891
rect 19681 845 19727 891
rect 19805 845 19851 891
rect 19929 845 19975 891
rect 20053 845 20099 891
rect 20177 845 20223 891
rect 20301 845 20347 891
rect 20425 845 20471 891
rect 20549 845 20595 891
rect 20673 845 20719 891
rect 20797 845 20843 891
rect 20921 845 20967 891
rect 21045 845 21091 891
rect 21169 845 21215 891
rect 21293 845 21339 891
rect 21417 845 21463 891
rect 21541 845 21587 891
rect 21665 845 21711 891
rect 21789 845 21835 891
rect 21913 845 21959 891
rect 22037 845 22083 891
rect 22161 845 22207 891
rect 22285 845 22331 891
rect 22409 845 22455 891
rect 22533 845 22579 891
rect 22657 845 22703 891
rect 22781 845 22827 891
rect 22905 845 22951 891
rect 23029 845 23075 891
rect 23153 845 23199 891
rect 23277 845 23323 891
rect 23401 845 23447 891
rect 23525 845 23571 891
rect 23649 845 23695 891
rect 23773 845 23819 891
rect 23897 845 23943 891
rect 24021 845 24067 891
rect 24145 845 24191 891
rect 24269 845 24315 891
rect 24393 845 24439 891
rect 24517 845 24563 891
rect 24641 845 24687 891
rect 24765 845 24811 891
rect 24889 845 24935 891
rect 25013 845 25059 891
rect 25137 845 25183 891
rect 25261 845 25307 891
rect 25385 845 25431 891
rect 25509 845 25555 891
rect 25633 845 25679 891
rect 25757 845 25803 891
rect 25881 845 25927 891
rect 26005 845 26051 891
rect 26129 845 26175 891
rect 26253 845 26299 891
rect 26377 845 26423 891
rect 26501 845 26547 891
rect 26625 845 26671 891
rect 26749 845 26795 891
rect 26873 845 26919 891
rect 26997 845 27043 891
rect 27121 845 27167 891
rect 27245 845 27291 891
rect 27369 845 27415 891
rect 27493 845 27539 891
rect 27617 845 27663 891
rect 27741 845 27787 891
rect 27865 845 27911 891
rect 27989 845 28035 891
rect 28113 845 28159 891
rect 28237 845 28283 891
rect 28361 845 28407 891
rect 28485 845 28531 891
rect 28609 845 28655 891
rect 28733 845 28779 891
rect 28857 845 28903 891
rect 28981 845 29027 891
rect 29105 845 29151 891
rect 29229 845 29275 891
rect 29353 845 29399 891
rect 29477 845 29523 891
rect 29601 845 29647 891
rect 29725 845 29771 891
rect 29849 845 29895 891
rect 29973 845 30019 891
rect 30097 845 30143 891
rect 30221 845 30267 891
rect 30345 845 30391 891
rect 30469 845 30515 891
rect 30593 845 30639 891
rect 30717 845 30763 891
rect 30841 845 30887 891
rect 30965 845 31011 891
rect 31089 845 31135 891
rect 31213 845 31259 891
rect 31337 845 31383 891
rect 31461 845 31507 891
rect 31585 845 31631 891
rect 31709 845 31755 891
rect 31833 845 31879 891
rect 31957 845 32003 891
rect 32081 845 32127 891
rect 32205 845 32251 891
rect 32329 845 32375 891
rect 32453 845 32499 891
rect 32577 845 32623 891
rect 32701 845 32747 891
rect 32825 845 32871 891
rect 32949 845 32995 891
rect 33073 845 33119 891
rect 33197 845 33243 891
rect 33321 845 33367 891
rect 33445 845 33491 891
rect 33569 845 33615 891
rect 33693 845 33739 891
rect 33817 845 33863 891
rect 33941 845 33987 891
rect 34065 845 34111 891
rect 34189 845 34235 891
rect 34313 845 34359 891
rect 34437 845 34483 891
rect 34561 845 34607 891
rect 34685 845 34731 891
rect 34809 845 34855 891
rect 34933 845 34979 891
rect 35057 845 35103 891
rect 35181 845 35227 891
rect 35305 845 35351 891
rect 35429 845 35475 891
rect 35553 845 35599 891
rect 35677 845 35723 891
rect 35801 845 35847 891
rect 35925 845 35971 891
rect 36049 845 36095 891
rect 36173 845 36219 891
rect 36297 845 36343 891
rect 36421 845 36467 891
rect 36545 845 36591 891
rect 36669 845 36715 891
rect 36793 845 36839 891
rect 36917 845 36963 891
rect 37041 845 37087 891
rect 37165 845 37211 891
rect 37289 845 37335 891
rect 37413 845 37459 891
rect 37537 845 37583 891
rect 37661 845 37707 891
rect 37785 845 37831 891
rect 37909 845 37955 891
rect 38033 845 38079 891
rect 38157 845 38203 891
rect 38281 845 38327 891
rect 38405 845 38451 891
rect 38529 845 38575 891
rect 38653 845 38699 891
rect 38777 845 38823 891
rect 38901 845 38947 891
rect 39025 845 39071 891
rect 39149 845 39195 891
rect 39273 845 39319 891
rect 39397 845 39443 891
rect 39521 845 39567 891
rect 39645 845 39691 891
rect 39769 845 39815 891
rect 39893 845 39939 891
rect 40017 845 40063 891
rect 40141 845 40187 891
rect 40265 845 40311 891
rect 40389 845 40435 891
rect 40513 845 40559 891
rect 40637 845 40683 891
rect 40761 845 40807 891
rect 40885 845 40931 891
rect 41009 845 41055 891
rect 41133 845 41179 891
rect 41257 845 41303 891
rect 41381 845 41427 891
rect 41505 845 41551 891
rect 41629 845 41675 891
rect 41753 845 41799 891
rect 41877 845 41923 891
rect 42001 845 42047 891
rect 42125 845 42171 891
rect 42249 845 42295 891
rect 42373 845 42419 891
rect 42497 845 42543 891
rect 42621 845 42667 891
rect 42745 845 42791 891
rect 42869 845 42915 891
rect 42993 845 43039 891
rect 43117 845 43163 891
rect 43241 845 43287 891
rect 43365 845 43411 891
rect 43489 845 43535 891
rect 43613 845 43659 891
rect 43737 845 43783 891
rect 43861 845 43907 891
rect 43985 845 44031 891
rect 44109 845 44155 891
rect 44233 845 44279 891
rect 44357 845 44403 891
rect 44481 845 44527 891
rect 44605 845 44651 891
rect 44729 845 44775 891
rect 44853 845 44899 891
rect 44977 845 45023 891
rect 45101 845 45147 891
rect 45225 845 45271 891
rect 45349 845 45395 891
rect 45473 845 45519 891
rect 45597 845 45643 891
rect 45721 845 45767 891
rect 45845 845 45891 891
rect 45969 845 46015 891
rect 46093 845 46139 891
rect 46217 845 46263 891
rect 46341 845 46387 891
rect 46465 845 46511 891
rect 46589 845 46635 891
rect 46713 845 46759 891
rect 46837 845 46883 891
rect 46961 845 47007 891
rect 47085 845 47131 891
rect 47209 845 47255 891
rect 47333 845 47379 891
rect 47457 845 47503 891
rect 47581 845 47627 891
rect 47705 845 47751 891
rect 47829 845 47875 891
rect 47953 845 47999 891
rect 48077 845 48123 891
rect 48201 845 48247 891
rect 48325 845 48371 891
rect 48449 845 48495 891
rect 48573 845 48619 891
rect 48697 845 48743 891
rect 48821 845 48867 891
rect 48945 845 48991 891
rect 49069 845 49115 891
rect 49193 845 49239 891
rect 49317 845 49363 891
rect 49441 845 49487 891
rect 49565 845 49611 891
rect 49689 845 49735 891
rect 49813 845 49859 891
rect 49937 845 49983 891
rect 50061 845 50107 891
rect 50185 845 50231 891
rect 50309 845 50355 891
rect 50433 845 50479 891
rect 50557 845 50603 891
rect 50681 845 50727 891
rect 50805 845 50851 891
rect 50929 845 50975 891
rect 51053 845 51099 891
rect 51177 845 51223 891
rect 51301 845 51347 891
rect 51425 845 51471 891
rect 51549 845 51595 891
rect 51673 845 51719 891
rect 51797 845 51843 891
rect 51921 845 51967 891
rect 52045 845 52091 891
rect 52169 845 52215 891
rect 52293 845 52339 891
rect 52417 845 52463 891
rect 52541 845 52587 891
rect 52665 845 52711 891
rect 52789 845 52835 891
rect 52913 845 52959 891
rect 53037 845 53083 891
rect 53161 845 53207 891
rect 53285 845 53331 891
rect 53409 845 53455 891
rect 53533 845 53579 891
rect 53657 845 53703 891
rect 53781 845 53827 891
rect 53905 845 53951 891
rect 54029 845 54075 891
rect 54153 845 54199 891
rect 54277 845 54323 891
rect 54401 845 54447 891
rect 54525 845 54571 891
rect 54649 845 54695 891
rect 54773 845 54819 891
rect 54897 845 54943 891
rect 55021 845 55067 891
rect 55145 845 55191 891
rect 55269 845 55315 891
rect 55393 845 55439 891
rect 55517 845 55563 891
rect 55641 845 55687 891
rect 55765 845 55811 891
rect 55889 845 55935 891
rect 56013 845 56059 891
rect 56137 845 56183 891
rect 56261 845 56307 891
rect 56385 845 56431 891
rect 56509 845 56555 891
rect 56633 845 56679 891
rect 56757 845 56803 891
rect 56881 845 56927 891
rect 57005 845 57051 891
rect 57129 845 57175 891
rect 57253 845 57299 891
rect 57377 845 57423 891
rect 57501 845 57547 891
rect 57625 845 57671 891
rect 57749 845 57795 891
rect 57873 845 57919 891
rect 57997 845 58043 891
rect 58121 845 58167 891
rect 58245 845 58291 891
rect 58369 845 58415 891
rect 58493 845 58539 891
rect 58617 845 58663 891
rect 58741 845 58787 891
rect 58865 845 58911 891
rect 58989 845 59035 891
rect 59113 845 59159 891
rect 59237 845 59283 891
rect 59361 845 59407 891
rect 59485 845 59531 891
rect 59609 845 59655 891
rect 59733 845 59779 891
rect 59857 845 59903 891
rect 59981 845 60027 891
rect 60105 845 60151 891
rect 60229 845 60275 891
rect 60353 845 60399 891
rect 60477 845 60523 891
rect 60601 845 60647 891
rect 60725 845 60771 891
rect 60849 845 60895 891
rect 60973 845 61019 891
rect 61097 845 61143 891
rect 61221 845 61267 891
rect 61345 845 61391 891
rect 61469 845 61515 891
rect 61593 845 61639 891
rect 61717 845 61763 891
rect 61841 845 61887 891
rect 61965 845 62011 891
rect 62089 845 62135 891
rect 62213 845 62259 891
rect 62337 845 62383 891
rect 62461 845 62507 891
rect 62585 845 62631 891
rect 62709 845 62755 891
rect 62833 845 62879 891
rect 62957 845 63003 891
rect 63081 845 63127 891
rect 63205 845 63251 891
rect 63329 845 63375 891
rect 63453 845 63499 891
rect 63577 845 63623 891
rect 63701 845 63747 891
rect 63825 845 63871 891
rect 63949 845 63995 891
rect 64073 845 64119 891
rect 64197 845 64243 891
rect 64321 845 64367 891
rect 64445 845 64491 891
rect 64569 845 64615 891
rect 64693 845 64739 891
rect 64817 845 64863 891
rect 64941 845 64987 891
rect 65065 845 65111 891
rect 65189 845 65235 891
rect 65313 845 65359 891
rect 65437 845 65483 891
rect 65561 845 65607 891
rect 65685 845 65731 891
rect 65809 845 65855 891
rect 65933 845 65979 891
rect 66057 845 66103 891
rect 66181 845 66227 891
rect 66305 845 66351 891
rect 66429 845 66475 891
rect 66553 845 66599 891
rect 66677 845 66723 891
rect 66801 845 66847 891
rect 66925 845 66971 891
rect 67049 845 67095 891
rect 67173 845 67219 891
rect 67297 845 67343 891
rect 67421 845 67467 891
rect 67545 845 67591 891
rect 67669 845 67715 891
rect 67793 845 67839 891
rect 67917 845 67963 891
rect 68041 845 68087 891
rect 68165 845 68211 891
rect 68289 845 68335 891
rect 68413 845 68459 891
rect 68537 845 68583 891
rect 68661 845 68707 891
rect 68785 845 68831 891
rect 68909 845 68955 891
rect 69033 845 69079 891
rect 69157 845 69203 891
rect 69281 845 69327 891
rect 69405 845 69451 891
rect 69529 845 69575 891
rect 69653 845 69699 891
rect 69777 845 69823 891
rect 69901 845 69947 891
rect 70025 845 70071 891
rect 70149 845 70195 891
rect 70273 845 70319 891
rect 70397 845 70443 891
rect 70521 845 70567 891
rect 70645 845 70691 891
rect 70769 845 70815 891
rect 70893 845 70939 891
rect 71017 845 71063 891
rect 71141 845 71187 891
rect 71265 845 71311 891
rect 71389 845 71435 891
rect 71513 845 71559 891
rect 71637 845 71683 891
rect 71761 845 71807 891
rect 71885 845 71931 891
rect 72009 845 72055 891
rect 72133 845 72179 891
rect 72257 845 72303 891
rect 72381 845 72427 891
rect 72505 845 72551 891
rect 72629 845 72675 891
rect 72753 845 72799 891
rect 72877 845 72923 891
rect 73001 845 73047 891
rect 73125 845 73171 891
rect 73249 845 73295 891
rect 73373 845 73419 891
rect 73497 845 73543 891
rect 73621 845 73667 891
rect 73745 845 73791 891
rect 73869 845 73915 891
rect 73993 845 74039 891
rect 74117 845 74163 891
rect 74241 845 74287 891
rect 74365 845 74411 891
rect 74489 845 74535 891
rect 74613 845 74659 891
rect 74737 845 74783 891
rect 74861 845 74907 891
rect 74985 845 75031 891
rect 75109 845 75155 891
rect 75233 845 75279 891
rect 75357 845 75403 891
rect 75481 845 75527 891
rect 75605 845 75651 891
rect 75729 845 75775 891
rect 75853 845 75899 891
rect 75977 845 76023 891
rect 76101 845 76147 891
rect 76225 845 76271 891
rect 76349 845 76395 891
rect 76473 845 76519 891
rect 76597 845 76643 891
rect 76721 845 76767 891
rect 76845 845 76891 891
rect 76969 845 77015 891
rect 77093 845 77139 891
rect 77217 845 77263 891
rect 77341 845 77387 891
rect 77465 845 77511 891
rect 77589 845 77635 891
rect 77713 845 77759 891
rect 77837 845 77883 891
rect 77961 845 78007 891
rect 78085 845 78131 891
rect 78209 845 78255 891
rect 78333 845 78379 891
rect 78457 845 78503 891
rect 78581 845 78627 891
rect 78705 845 78751 891
rect 78829 845 78875 891
rect 78953 845 78999 891
rect 79077 845 79123 891
rect 79201 845 79247 891
rect 79325 845 79371 891
rect 79449 845 79495 891
rect 79573 845 79619 891
rect 79697 845 79743 891
rect 79821 845 79867 891
rect 79945 845 79991 891
rect 80069 845 80115 891
rect 80193 845 80239 891
rect 80317 845 80363 891
rect 80441 845 80487 891
rect 80565 845 80611 891
rect 80689 845 80735 891
rect 80813 845 80859 891
rect 80937 845 80983 891
rect 81061 845 81107 891
rect 81185 845 81231 891
rect 81309 845 81355 891
rect 81433 845 81479 891
rect 81557 845 81603 891
rect 81681 845 81727 891
rect 81805 845 81851 891
rect 81929 845 81975 891
rect 82053 845 82099 891
rect 82177 845 82223 891
rect 82301 845 82347 891
rect 82425 845 82471 891
rect 82549 845 82595 891
rect 82673 845 82719 891
rect 82797 845 82843 891
rect 82921 845 82967 891
rect 83045 845 83091 891
rect 83169 845 83215 891
rect 83293 845 83339 891
rect 83417 845 83463 891
rect 83541 845 83587 891
rect 83665 845 83711 891
rect 83789 845 83835 891
rect 83913 845 83959 891
rect 84037 845 84083 891
rect 84161 845 84207 891
rect 84285 845 84331 891
rect 84409 845 84455 891
rect 84533 845 84579 891
rect 84657 845 84703 891
rect 84781 845 84827 891
rect 84905 845 84951 891
rect 85029 845 85075 891
rect 85153 845 85199 891
rect 85277 845 85323 891
rect 85401 845 85447 891
rect 85525 845 85571 891
rect 85649 845 85695 891
rect 89 721 135 767
rect 213 721 259 767
rect 337 721 383 767
rect 461 721 507 767
rect 585 721 631 767
rect 709 721 755 767
rect 833 721 879 767
rect 957 721 1003 767
rect 1081 721 1127 767
rect 1205 721 1251 767
rect 1329 721 1375 767
rect 1453 721 1499 767
rect 1577 721 1623 767
rect 1701 721 1747 767
rect 1825 721 1871 767
rect 1949 721 1995 767
rect 2073 721 2119 767
rect 2197 721 2243 767
rect 2321 721 2367 767
rect 2445 721 2491 767
rect 2569 721 2615 767
rect 2693 721 2739 767
rect 2817 721 2863 767
rect 2941 721 2987 767
rect 3065 721 3111 767
rect 3189 721 3235 767
rect 3313 721 3359 767
rect 3437 721 3483 767
rect 3561 721 3607 767
rect 3685 721 3731 767
rect 3809 721 3855 767
rect 3933 721 3979 767
rect 4057 721 4103 767
rect 4181 721 4227 767
rect 4305 721 4351 767
rect 4429 721 4475 767
rect 4553 721 4599 767
rect 4677 721 4723 767
rect 4801 721 4847 767
rect 4925 721 4971 767
rect 5049 721 5095 767
rect 5173 721 5219 767
rect 5297 721 5343 767
rect 5421 721 5467 767
rect 5545 721 5591 767
rect 5669 721 5715 767
rect 5793 721 5839 767
rect 5917 721 5963 767
rect 6041 721 6087 767
rect 6165 721 6211 767
rect 6289 721 6335 767
rect 6413 721 6459 767
rect 6537 721 6583 767
rect 6661 721 6707 767
rect 6785 721 6831 767
rect 6909 721 6955 767
rect 7033 721 7079 767
rect 7157 721 7203 767
rect 7281 721 7327 767
rect 7405 721 7451 767
rect 7529 721 7575 767
rect 7653 721 7699 767
rect 7777 721 7823 767
rect 7901 721 7947 767
rect 8025 721 8071 767
rect 8149 721 8195 767
rect 8273 721 8319 767
rect 8397 721 8443 767
rect 8521 721 8567 767
rect 8645 721 8691 767
rect 8769 721 8815 767
rect 8893 721 8939 767
rect 9017 721 9063 767
rect 9141 721 9187 767
rect 9265 721 9311 767
rect 9389 721 9435 767
rect 9513 721 9559 767
rect 9637 721 9683 767
rect 9761 721 9807 767
rect 9885 721 9931 767
rect 10009 721 10055 767
rect 10133 721 10179 767
rect 10257 721 10303 767
rect 10381 721 10427 767
rect 10505 721 10551 767
rect 10629 721 10675 767
rect 10753 721 10799 767
rect 10877 721 10923 767
rect 11001 721 11047 767
rect 11125 721 11171 767
rect 11249 721 11295 767
rect 11373 721 11419 767
rect 11497 721 11543 767
rect 11621 721 11667 767
rect 11745 721 11791 767
rect 11869 721 11915 767
rect 11993 721 12039 767
rect 12117 721 12163 767
rect 12241 721 12287 767
rect 12365 721 12411 767
rect 12489 721 12535 767
rect 12613 721 12659 767
rect 12737 721 12783 767
rect 12861 721 12907 767
rect 12985 721 13031 767
rect 13109 721 13155 767
rect 13233 721 13279 767
rect 13357 721 13403 767
rect 13481 721 13527 767
rect 13605 721 13651 767
rect 13729 721 13775 767
rect 13853 721 13899 767
rect 13977 721 14023 767
rect 14101 721 14147 767
rect 14225 721 14271 767
rect 14349 721 14395 767
rect 14473 721 14519 767
rect 14597 721 14643 767
rect 14721 721 14767 767
rect 14845 721 14891 767
rect 14969 721 15015 767
rect 15093 721 15139 767
rect 15217 721 15263 767
rect 15341 721 15387 767
rect 15465 721 15511 767
rect 15589 721 15635 767
rect 15713 721 15759 767
rect 15837 721 15883 767
rect 15961 721 16007 767
rect 16085 721 16131 767
rect 16209 721 16255 767
rect 16333 721 16379 767
rect 16457 721 16503 767
rect 16581 721 16627 767
rect 16705 721 16751 767
rect 16829 721 16875 767
rect 16953 721 16999 767
rect 17077 721 17123 767
rect 17201 721 17247 767
rect 17325 721 17371 767
rect 17449 721 17495 767
rect 17573 721 17619 767
rect 17697 721 17743 767
rect 17821 721 17867 767
rect 17945 721 17991 767
rect 18069 721 18115 767
rect 18193 721 18239 767
rect 18317 721 18363 767
rect 18441 721 18487 767
rect 18565 721 18611 767
rect 18689 721 18735 767
rect 18813 721 18859 767
rect 18937 721 18983 767
rect 19061 721 19107 767
rect 19185 721 19231 767
rect 19309 721 19355 767
rect 19433 721 19479 767
rect 19557 721 19603 767
rect 19681 721 19727 767
rect 19805 721 19851 767
rect 19929 721 19975 767
rect 20053 721 20099 767
rect 20177 721 20223 767
rect 20301 721 20347 767
rect 20425 721 20471 767
rect 20549 721 20595 767
rect 20673 721 20719 767
rect 20797 721 20843 767
rect 20921 721 20967 767
rect 21045 721 21091 767
rect 21169 721 21215 767
rect 21293 721 21339 767
rect 21417 721 21463 767
rect 21541 721 21587 767
rect 21665 721 21711 767
rect 21789 721 21835 767
rect 21913 721 21959 767
rect 22037 721 22083 767
rect 22161 721 22207 767
rect 22285 721 22331 767
rect 22409 721 22455 767
rect 22533 721 22579 767
rect 22657 721 22703 767
rect 22781 721 22827 767
rect 22905 721 22951 767
rect 23029 721 23075 767
rect 23153 721 23199 767
rect 23277 721 23323 767
rect 23401 721 23447 767
rect 23525 721 23571 767
rect 23649 721 23695 767
rect 23773 721 23819 767
rect 23897 721 23943 767
rect 24021 721 24067 767
rect 24145 721 24191 767
rect 24269 721 24315 767
rect 24393 721 24439 767
rect 24517 721 24563 767
rect 24641 721 24687 767
rect 24765 721 24811 767
rect 24889 721 24935 767
rect 25013 721 25059 767
rect 25137 721 25183 767
rect 25261 721 25307 767
rect 25385 721 25431 767
rect 25509 721 25555 767
rect 25633 721 25679 767
rect 25757 721 25803 767
rect 25881 721 25927 767
rect 26005 721 26051 767
rect 26129 721 26175 767
rect 26253 721 26299 767
rect 26377 721 26423 767
rect 26501 721 26547 767
rect 26625 721 26671 767
rect 26749 721 26795 767
rect 26873 721 26919 767
rect 26997 721 27043 767
rect 27121 721 27167 767
rect 27245 721 27291 767
rect 27369 721 27415 767
rect 27493 721 27539 767
rect 27617 721 27663 767
rect 27741 721 27787 767
rect 27865 721 27911 767
rect 27989 721 28035 767
rect 28113 721 28159 767
rect 28237 721 28283 767
rect 28361 721 28407 767
rect 28485 721 28531 767
rect 28609 721 28655 767
rect 28733 721 28779 767
rect 28857 721 28903 767
rect 28981 721 29027 767
rect 29105 721 29151 767
rect 29229 721 29275 767
rect 29353 721 29399 767
rect 29477 721 29523 767
rect 29601 721 29647 767
rect 29725 721 29771 767
rect 29849 721 29895 767
rect 29973 721 30019 767
rect 30097 721 30143 767
rect 30221 721 30267 767
rect 30345 721 30391 767
rect 30469 721 30515 767
rect 30593 721 30639 767
rect 30717 721 30763 767
rect 30841 721 30887 767
rect 30965 721 31011 767
rect 31089 721 31135 767
rect 31213 721 31259 767
rect 31337 721 31383 767
rect 31461 721 31507 767
rect 31585 721 31631 767
rect 31709 721 31755 767
rect 31833 721 31879 767
rect 31957 721 32003 767
rect 32081 721 32127 767
rect 32205 721 32251 767
rect 32329 721 32375 767
rect 32453 721 32499 767
rect 32577 721 32623 767
rect 32701 721 32747 767
rect 32825 721 32871 767
rect 32949 721 32995 767
rect 33073 721 33119 767
rect 33197 721 33243 767
rect 33321 721 33367 767
rect 33445 721 33491 767
rect 33569 721 33615 767
rect 33693 721 33739 767
rect 33817 721 33863 767
rect 33941 721 33987 767
rect 34065 721 34111 767
rect 34189 721 34235 767
rect 34313 721 34359 767
rect 34437 721 34483 767
rect 34561 721 34607 767
rect 34685 721 34731 767
rect 34809 721 34855 767
rect 34933 721 34979 767
rect 35057 721 35103 767
rect 35181 721 35227 767
rect 35305 721 35351 767
rect 35429 721 35475 767
rect 35553 721 35599 767
rect 35677 721 35723 767
rect 35801 721 35847 767
rect 35925 721 35971 767
rect 36049 721 36095 767
rect 36173 721 36219 767
rect 36297 721 36343 767
rect 36421 721 36467 767
rect 36545 721 36591 767
rect 36669 721 36715 767
rect 36793 721 36839 767
rect 36917 721 36963 767
rect 37041 721 37087 767
rect 37165 721 37211 767
rect 37289 721 37335 767
rect 37413 721 37459 767
rect 37537 721 37583 767
rect 37661 721 37707 767
rect 37785 721 37831 767
rect 37909 721 37955 767
rect 38033 721 38079 767
rect 38157 721 38203 767
rect 38281 721 38327 767
rect 38405 721 38451 767
rect 38529 721 38575 767
rect 38653 721 38699 767
rect 38777 721 38823 767
rect 38901 721 38947 767
rect 39025 721 39071 767
rect 39149 721 39195 767
rect 39273 721 39319 767
rect 39397 721 39443 767
rect 39521 721 39567 767
rect 39645 721 39691 767
rect 39769 721 39815 767
rect 39893 721 39939 767
rect 40017 721 40063 767
rect 40141 721 40187 767
rect 40265 721 40311 767
rect 40389 721 40435 767
rect 40513 721 40559 767
rect 40637 721 40683 767
rect 40761 721 40807 767
rect 40885 721 40931 767
rect 41009 721 41055 767
rect 41133 721 41179 767
rect 41257 721 41303 767
rect 41381 721 41427 767
rect 41505 721 41551 767
rect 41629 721 41675 767
rect 41753 721 41799 767
rect 41877 721 41923 767
rect 42001 721 42047 767
rect 42125 721 42171 767
rect 42249 721 42295 767
rect 42373 721 42419 767
rect 42497 721 42543 767
rect 42621 721 42667 767
rect 42745 721 42791 767
rect 42869 721 42915 767
rect 42993 721 43039 767
rect 43117 721 43163 767
rect 43241 721 43287 767
rect 43365 721 43411 767
rect 43489 721 43535 767
rect 43613 721 43659 767
rect 43737 721 43783 767
rect 43861 721 43907 767
rect 43985 721 44031 767
rect 44109 721 44155 767
rect 44233 721 44279 767
rect 44357 721 44403 767
rect 44481 721 44527 767
rect 44605 721 44651 767
rect 44729 721 44775 767
rect 44853 721 44899 767
rect 44977 721 45023 767
rect 45101 721 45147 767
rect 45225 721 45271 767
rect 45349 721 45395 767
rect 45473 721 45519 767
rect 45597 721 45643 767
rect 45721 721 45767 767
rect 45845 721 45891 767
rect 45969 721 46015 767
rect 46093 721 46139 767
rect 46217 721 46263 767
rect 46341 721 46387 767
rect 46465 721 46511 767
rect 46589 721 46635 767
rect 46713 721 46759 767
rect 46837 721 46883 767
rect 46961 721 47007 767
rect 47085 721 47131 767
rect 47209 721 47255 767
rect 47333 721 47379 767
rect 47457 721 47503 767
rect 47581 721 47627 767
rect 47705 721 47751 767
rect 47829 721 47875 767
rect 47953 721 47999 767
rect 48077 721 48123 767
rect 48201 721 48247 767
rect 48325 721 48371 767
rect 48449 721 48495 767
rect 48573 721 48619 767
rect 48697 721 48743 767
rect 48821 721 48867 767
rect 48945 721 48991 767
rect 49069 721 49115 767
rect 49193 721 49239 767
rect 49317 721 49363 767
rect 49441 721 49487 767
rect 49565 721 49611 767
rect 49689 721 49735 767
rect 49813 721 49859 767
rect 49937 721 49983 767
rect 50061 721 50107 767
rect 50185 721 50231 767
rect 50309 721 50355 767
rect 50433 721 50479 767
rect 50557 721 50603 767
rect 50681 721 50727 767
rect 50805 721 50851 767
rect 50929 721 50975 767
rect 51053 721 51099 767
rect 51177 721 51223 767
rect 51301 721 51347 767
rect 51425 721 51471 767
rect 51549 721 51595 767
rect 51673 721 51719 767
rect 51797 721 51843 767
rect 51921 721 51967 767
rect 52045 721 52091 767
rect 52169 721 52215 767
rect 52293 721 52339 767
rect 52417 721 52463 767
rect 52541 721 52587 767
rect 52665 721 52711 767
rect 52789 721 52835 767
rect 52913 721 52959 767
rect 53037 721 53083 767
rect 53161 721 53207 767
rect 53285 721 53331 767
rect 53409 721 53455 767
rect 53533 721 53579 767
rect 53657 721 53703 767
rect 53781 721 53827 767
rect 53905 721 53951 767
rect 54029 721 54075 767
rect 54153 721 54199 767
rect 54277 721 54323 767
rect 54401 721 54447 767
rect 54525 721 54571 767
rect 54649 721 54695 767
rect 54773 721 54819 767
rect 54897 721 54943 767
rect 55021 721 55067 767
rect 55145 721 55191 767
rect 55269 721 55315 767
rect 55393 721 55439 767
rect 55517 721 55563 767
rect 55641 721 55687 767
rect 55765 721 55811 767
rect 55889 721 55935 767
rect 56013 721 56059 767
rect 56137 721 56183 767
rect 56261 721 56307 767
rect 56385 721 56431 767
rect 56509 721 56555 767
rect 56633 721 56679 767
rect 56757 721 56803 767
rect 56881 721 56927 767
rect 57005 721 57051 767
rect 57129 721 57175 767
rect 57253 721 57299 767
rect 57377 721 57423 767
rect 57501 721 57547 767
rect 57625 721 57671 767
rect 57749 721 57795 767
rect 57873 721 57919 767
rect 57997 721 58043 767
rect 58121 721 58167 767
rect 58245 721 58291 767
rect 58369 721 58415 767
rect 58493 721 58539 767
rect 58617 721 58663 767
rect 58741 721 58787 767
rect 58865 721 58911 767
rect 58989 721 59035 767
rect 59113 721 59159 767
rect 59237 721 59283 767
rect 59361 721 59407 767
rect 59485 721 59531 767
rect 59609 721 59655 767
rect 59733 721 59779 767
rect 59857 721 59903 767
rect 59981 721 60027 767
rect 60105 721 60151 767
rect 60229 721 60275 767
rect 60353 721 60399 767
rect 60477 721 60523 767
rect 60601 721 60647 767
rect 60725 721 60771 767
rect 60849 721 60895 767
rect 60973 721 61019 767
rect 61097 721 61143 767
rect 61221 721 61267 767
rect 61345 721 61391 767
rect 61469 721 61515 767
rect 61593 721 61639 767
rect 61717 721 61763 767
rect 61841 721 61887 767
rect 61965 721 62011 767
rect 62089 721 62135 767
rect 62213 721 62259 767
rect 62337 721 62383 767
rect 62461 721 62507 767
rect 62585 721 62631 767
rect 62709 721 62755 767
rect 62833 721 62879 767
rect 62957 721 63003 767
rect 63081 721 63127 767
rect 63205 721 63251 767
rect 63329 721 63375 767
rect 63453 721 63499 767
rect 63577 721 63623 767
rect 63701 721 63747 767
rect 63825 721 63871 767
rect 63949 721 63995 767
rect 64073 721 64119 767
rect 64197 721 64243 767
rect 64321 721 64367 767
rect 64445 721 64491 767
rect 64569 721 64615 767
rect 64693 721 64739 767
rect 64817 721 64863 767
rect 64941 721 64987 767
rect 65065 721 65111 767
rect 65189 721 65235 767
rect 65313 721 65359 767
rect 65437 721 65483 767
rect 65561 721 65607 767
rect 65685 721 65731 767
rect 65809 721 65855 767
rect 65933 721 65979 767
rect 66057 721 66103 767
rect 66181 721 66227 767
rect 66305 721 66351 767
rect 66429 721 66475 767
rect 66553 721 66599 767
rect 66677 721 66723 767
rect 66801 721 66847 767
rect 66925 721 66971 767
rect 67049 721 67095 767
rect 67173 721 67219 767
rect 67297 721 67343 767
rect 67421 721 67467 767
rect 67545 721 67591 767
rect 67669 721 67715 767
rect 67793 721 67839 767
rect 67917 721 67963 767
rect 68041 721 68087 767
rect 68165 721 68211 767
rect 68289 721 68335 767
rect 68413 721 68459 767
rect 68537 721 68583 767
rect 68661 721 68707 767
rect 68785 721 68831 767
rect 68909 721 68955 767
rect 69033 721 69079 767
rect 69157 721 69203 767
rect 69281 721 69327 767
rect 69405 721 69451 767
rect 69529 721 69575 767
rect 69653 721 69699 767
rect 69777 721 69823 767
rect 69901 721 69947 767
rect 70025 721 70071 767
rect 70149 721 70195 767
rect 70273 721 70319 767
rect 70397 721 70443 767
rect 70521 721 70567 767
rect 70645 721 70691 767
rect 70769 721 70815 767
rect 70893 721 70939 767
rect 71017 721 71063 767
rect 71141 721 71187 767
rect 71265 721 71311 767
rect 71389 721 71435 767
rect 71513 721 71559 767
rect 71637 721 71683 767
rect 71761 721 71807 767
rect 71885 721 71931 767
rect 72009 721 72055 767
rect 72133 721 72179 767
rect 72257 721 72303 767
rect 72381 721 72427 767
rect 72505 721 72551 767
rect 72629 721 72675 767
rect 72753 721 72799 767
rect 72877 721 72923 767
rect 73001 721 73047 767
rect 73125 721 73171 767
rect 73249 721 73295 767
rect 73373 721 73419 767
rect 73497 721 73543 767
rect 73621 721 73667 767
rect 73745 721 73791 767
rect 73869 721 73915 767
rect 73993 721 74039 767
rect 74117 721 74163 767
rect 74241 721 74287 767
rect 74365 721 74411 767
rect 74489 721 74535 767
rect 74613 721 74659 767
rect 74737 721 74783 767
rect 74861 721 74907 767
rect 74985 721 75031 767
rect 75109 721 75155 767
rect 75233 721 75279 767
rect 75357 721 75403 767
rect 75481 721 75527 767
rect 75605 721 75651 767
rect 75729 721 75775 767
rect 75853 721 75899 767
rect 75977 721 76023 767
rect 76101 721 76147 767
rect 76225 721 76271 767
rect 76349 721 76395 767
rect 76473 721 76519 767
rect 76597 721 76643 767
rect 76721 721 76767 767
rect 76845 721 76891 767
rect 76969 721 77015 767
rect 77093 721 77139 767
rect 77217 721 77263 767
rect 77341 721 77387 767
rect 77465 721 77511 767
rect 77589 721 77635 767
rect 77713 721 77759 767
rect 77837 721 77883 767
rect 77961 721 78007 767
rect 78085 721 78131 767
rect 78209 721 78255 767
rect 78333 721 78379 767
rect 78457 721 78503 767
rect 78581 721 78627 767
rect 78705 721 78751 767
rect 78829 721 78875 767
rect 78953 721 78999 767
rect 79077 721 79123 767
rect 79201 721 79247 767
rect 79325 721 79371 767
rect 79449 721 79495 767
rect 79573 721 79619 767
rect 79697 721 79743 767
rect 79821 721 79867 767
rect 79945 721 79991 767
rect 80069 721 80115 767
rect 80193 721 80239 767
rect 80317 721 80363 767
rect 80441 721 80487 767
rect 80565 721 80611 767
rect 80689 721 80735 767
rect 80813 721 80859 767
rect 80937 721 80983 767
rect 81061 721 81107 767
rect 81185 721 81231 767
rect 81309 721 81355 767
rect 81433 721 81479 767
rect 81557 721 81603 767
rect 81681 721 81727 767
rect 81805 721 81851 767
rect 81929 721 81975 767
rect 82053 721 82099 767
rect 82177 721 82223 767
rect 82301 721 82347 767
rect 82425 721 82471 767
rect 82549 721 82595 767
rect 82673 721 82719 767
rect 82797 721 82843 767
rect 82921 721 82967 767
rect 83045 721 83091 767
rect 83169 721 83215 767
rect 83293 721 83339 767
rect 83417 721 83463 767
rect 83541 721 83587 767
rect 83665 721 83711 767
rect 83789 721 83835 767
rect 83913 721 83959 767
rect 84037 721 84083 767
rect 84161 721 84207 767
rect 84285 721 84331 767
rect 84409 721 84455 767
rect 84533 721 84579 767
rect 84657 721 84703 767
rect 84781 721 84827 767
rect 84905 721 84951 767
rect 85029 721 85075 767
rect 85153 721 85199 767
rect 85277 721 85323 767
rect 85401 721 85447 767
rect 85525 721 85571 767
rect 85649 721 85695 767
rect 89 597 135 643
rect 213 597 259 643
rect 337 597 383 643
rect 461 597 507 643
rect 585 597 631 643
rect 709 597 755 643
rect 833 597 879 643
rect 957 597 1003 643
rect 1081 597 1127 643
rect 1205 597 1251 643
rect 1329 597 1375 643
rect 1453 597 1499 643
rect 1577 597 1623 643
rect 1701 597 1747 643
rect 1825 597 1871 643
rect 1949 597 1995 643
rect 2073 597 2119 643
rect 2197 597 2243 643
rect 2321 597 2367 643
rect 2445 597 2491 643
rect 2569 597 2615 643
rect 2693 597 2739 643
rect 2817 597 2863 643
rect 2941 597 2987 643
rect 3065 597 3111 643
rect 3189 597 3235 643
rect 3313 597 3359 643
rect 3437 597 3483 643
rect 3561 597 3607 643
rect 3685 597 3731 643
rect 3809 597 3855 643
rect 3933 597 3979 643
rect 4057 597 4103 643
rect 4181 597 4227 643
rect 4305 597 4351 643
rect 4429 597 4475 643
rect 4553 597 4599 643
rect 4677 597 4723 643
rect 4801 597 4847 643
rect 4925 597 4971 643
rect 5049 597 5095 643
rect 5173 597 5219 643
rect 5297 597 5343 643
rect 5421 597 5467 643
rect 5545 597 5591 643
rect 5669 597 5715 643
rect 5793 597 5839 643
rect 5917 597 5963 643
rect 6041 597 6087 643
rect 6165 597 6211 643
rect 6289 597 6335 643
rect 6413 597 6459 643
rect 6537 597 6583 643
rect 6661 597 6707 643
rect 6785 597 6831 643
rect 6909 597 6955 643
rect 7033 597 7079 643
rect 7157 597 7203 643
rect 7281 597 7327 643
rect 7405 597 7451 643
rect 7529 597 7575 643
rect 7653 597 7699 643
rect 7777 597 7823 643
rect 7901 597 7947 643
rect 8025 597 8071 643
rect 8149 597 8195 643
rect 8273 597 8319 643
rect 8397 597 8443 643
rect 8521 597 8567 643
rect 8645 597 8691 643
rect 8769 597 8815 643
rect 8893 597 8939 643
rect 9017 597 9063 643
rect 9141 597 9187 643
rect 9265 597 9311 643
rect 9389 597 9435 643
rect 9513 597 9559 643
rect 9637 597 9683 643
rect 9761 597 9807 643
rect 9885 597 9931 643
rect 10009 597 10055 643
rect 10133 597 10179 643
rect 10257 597 10303 643
rect 10381 597 10427 643
rect 10505 597 10551 643
rect 10629 597 10675 643
rect 10753 597 10799 643
rect 10877 597 10923 643
rect 11001 597 11047 643
rect 11125 597 11171 643
rect 11249 597 11295 643
rect 11373 597 11419 643
rect 11497 597 11543 643
rect 11621 597 11667 643
rect 11745 597 11791 643
rect 11869 597 11915 643
rect 11993 597 12039 643
rect 12117 597 12163 643
rect 12241 597 12287 643
rect 12365 597 12411 643
rect 12489 597 12535 643
rect 12613 597 12659 643
rect 12737 597 12783 643
rect 12861 597 12907 643
rect 12985 597 13031 643
rect 13109 597 13155 643
rect 13233 597 13279 643
rect 13357 597 13403 643
rect 13481 597 13527 643
rect 13605 597 13651 643
rect 13729 597 13775 643
rect 13853 597 13899 643
rect 13977 597 14023 643
rect 14101 597 14147 643
rect 14225 597 14271 643
rect 14349 597 14395 643
rect 14473 597 14519 643
rect 14597 597 14643 643
rect 14721 597 14767 643
rect 14845 597 14891 643
rect 14969 597 15015 643
rect 15093 597 15139 643
rect 15217 597 15263 643
rect 15341 597 15387 643
rect 15465 597 15511 643
rect 15589 597 15635 643
rect 15713 597 15759 643
rect 15837 597 15883 643
rect 15961 597 16007 643
rect 16085 597 16131 643
rect 16209 597 16255 643
rect 16333 597 16379 643
rect 16457 597 16503 643
rect 16581 597 16627 643
rect 16705 597 16751 643
rect 16829 597 16875 643
rect 16953 597 16999 643
rect 17077 597 17123 643
rect 17201 597 17247 643
rect 17325 597 17371 643
rect 17449 597 17495 643
rect 17573 597 17619 643
rect 17697 597 17743 643
rect 17821 597 17867 643
rect 17945 597 17991 643
rect 18069 597 18115 643
rect 18193 597 18239 643
rect 18317 597 18363 643
rect 18441 597 18487 643
rect 18565 597 18611 643
rect 18689 597 18735 643
rect 18813 597 18859 643
rect 18937 597 18983 643
rect 19061 597 19107 643
rect 19185 597 19231 643
rect 19309 597 19355 643
rect 19433 597 19479 643
rect 19557 597 19603 643
rect 19681 597 19727 643
rect 19805 597 19851 643
rect 19929 597 19975 643
rect 20053 597 20099 643
rect 20177 597 20223 643
rect 20301 597 20347 643
rect 20425 597 20471 643
rect 20549 597 20595 643
rect 20673 597 20719 643
rect 20797 597 20843 643
rect 20921 597 20967 643
rect 21045 597 21091 643
rect 21169 597 21215 643
rect 21293 597 21339 643
rect 21417 597 21463 643
rect 21541 597 21587 643
rect 21665 597 21711 643
rect 21789 597 21835 643
rect 21913 597 21959 643
rect 22037 597 22083 643
rect 22161 597 22207 643
rect 22285 597 22331 643
rect 22409 597 22455 643
rect 22533 597 22579 643
rect 22657 597 22703 643
rect 22781 597 22827 643
rect 22905 597 22951 643
rect 23029 597 23075 643
rect 23153 597 23199 643
rect 23277 597 23323 643
rect 23401 597 23447 643
rect 23525 597 23571 643
rect 23649 597 23695 643
rect 23773 597 23819 643
rect 23897 597 23943 643
rect 24021 597 24067 643
rect 24145 597 24191 643
rect 24269 597 24315 643
rect 24393 597 24439 643
rect 24517 597 24563 643
rect 24641 597 24687 643
rect 24765 597 24811 643
rect 24889 597 24935 643
rect 25013 597 25059 643
rect 25137 597 25183 643
rect 25261 597 25307 643
rect 25385 597 25431 643
rect 25509 597 25555 643
rect 25633 597 25679 643
rect 25757 597 25803 643
rect 25881 597 25927 643
rect 26005 597 26051 643
rect 26129 597 26175 643
rect 26253 597 26299 643
rect 26377 597 26423 643
rect 26501 597 26547 643
rect 26625 597 26671 643
rect 26749 597 26795 643
rect 26873 597 26919 643
rect 26997 597 27043 643
rect 27121 597 27167 643
rect 27245 597 27291 643
rect 27369 597 27415 643
rect 27493 597 27539 643
rect 27617 597 27663 643
rect 27741 597 27787 643
rect 27865 597 27911 643
rect 27989 597 28035 643
rect 28113 597 28159 643
rect 28237 597 28283 643
rect 28361 597 28407 643
rect 28485 597 28531 643
rect 28609 597 28655 643
rect 28733 597 28779 643
rect 28857 597 28903 643
rect 28981 597 29027 643
rect 29105 597 29151 643
rect 29229 597 29275 643
rect 29353 597 29399 643
rect 29477 597 29523 643
rect 29601 597 29647 643
rect 29725 597 29771 643
rect 29849 597 29895 643
rect 29973 597 30019 643
rect 30097 597 30143 643
rect 30221 597 30267 643
rect 30345 597 30391 643
rect 30469 597 30515 643
rect 30593 597 30639 643
rect 30717 597 30763 643
rect 30841 597 30887 643
rect 30965 597 31011 643
rect 31089 597 31135 643
rect 31213 597 31259 643
rect 31337 597 31383 643
rect 31461 597 31507 643
rect 31585 597 31631 643
rect 31709 597 31755 643
rect 31833 597 31879 643
rect 31957 597 32003 643
rect 32081 597 32127 643
rect 32205 597 32251 643
rect 32329 597 32375 643
rect 32453 597 32499 643
rect 32577 597 32623 643
rect 32701 597 32747 643
rect 32825 597 32871 643
rect 32949 597 32995 643
rect 33073 597 33119 643
rect 33197 597 33243 643
rect 33321 597 33367 643
rect 33445 597 33491 643
rect 33569 597 33615 643
rect 33693 597 33739 643
rect 33817 597 33863 643
rect 33941 597 33987 643
rect 34065 597 34111 643
rect 34189 597 34235 643
rect 34313 597 34359 643
rect 34437 597 34483 643
rect 34561 597 34607 643
rect 34685 597 34731 643
rect 34809 597 34855 643
rect 34933 597 34979 643
rect 35057 597 35103 643
rect 35181 597 35227 643
rect 35305 597 35351 643
rect 35429 597 35475 643
rect 35553 597 35599 643
rect 35677 597 35723 643
rect 35801 597 35847 643
rect 35925 597 35971 643
rect 36049 597 36095 643
rect 36173 597 36219 643
rect 36297 597 36343 643
rect 36421 597 36467 643
rect 36545 597 36591 643
rect 36669 597 36715 643
rect 36793 597 36839 643
rect 36917 597 36963 643
rect 37041 597 37087 643
rect 37165 597 37211 643
rect 37289 597 37335 643
rect 37413 597 37459 643
rect 37537 597 37583 643
rect 37661 597 37707 643
rect 37785 597 37831 643
rect 37909 597 37955 643
rect 38033 597 38079 643
rect 38157 597 38203 643
rect 38281 597 38327 643
rect 38405 597 38451 643
rect 38529 597 38575 643
rect 38653 597 38699 643
rect 38777 597 38823 643
rect 38901 597 38947 643
rect 39025 597 39071 643
rect 39149 597 39195 643
rect 39273 597 39319 643
rect 39397 597 39443 643
rect 39521 597 39567 643
rect 39645 597 39691 643
rect 39769 597 39815 643
rect 39893 597 39939 643
rect 40017 597 40063 643
rect 40141 597 40187 643
rect 40265 597 40311 643
rect 40389 597 40435 643
rect 40513 597 40559 643
rect 40637 597 40683 643
rect 40761 597 40807 643
rect 40885 597 40931 643
rect 41009 597 41055 643
rect 41133 597 41179 643
rect 41257 597 41303 643
rect 41381 597 41427 643
rect 41505 597 41551 643
rect 41629 597 41675 643
rect 41753 597 41799 643
rect 41877 597 41923 643
rect 42001 597 42047 643
rect 42125 597 42171 643
rect 42249 597 42295 643
rect 42373 597 42419 643
rect 42497 597 42543 643
rect 42621 597 42667 643
rect 42745 597 42791 643
rect 42869 597 42915 643
rect 42993 597 43039 643
rect 43117 597 43163 643
rect 43241 597 43287 643
rect 43365 597 43411 643
rect 43489 597 43535 643
rect 43613 597 43659 643
rect 43737 597 43783 643
rect 43861 597 43907 643
rect 43985 597 44031 643
rect 44109 597 44155 643
rect 44233 597 44279 643
rect 44357 597 44403 643
rect 44481 597 44527 643
rect 44605 597 44651 643
rect 44729 597 44775 643
rect 44853 597 44899 643
rect 44977 597 45023 643
rect 45101 597 45147 643
rect 45225 597 45271 643
rect 45349 597 45395 643
rect 45473 597 45519 643
rect 45597 597 45643 643
rect 45721 597 45767 643
rect 45845 597 45891 643
rect 45969 597 46015 643
rect 46093 597 46139 643
rect 46217 597 46263 643
rect 46341 597 46387 643
rect 46465 597 46511 643
rect 46589 597 46635 643
rect 46713 597 46759 643
rect 46837 597 46883 643
rect 46961 597 47007 643
rect 47085 597 47131 643
rect 47209 597 47255 643
rect 47333 597 47379 643
rect 47457 597 47503 643
rect 47581 597 47627 643
rect 47705 597 47751 643
rect 47829 597 47875 643
rect 47953 597 47999 643
rect 48077 597 48123 643
rect 48201 597 48247 643
rect 48325 597 48371 643
rect 48449 597 48495 643
rect 48573 597 48619 643
rect 48697 597 48743 643
rect 48821 597 48867 643
rect 48945 597 48991 643
rect 49069 597 49115 643
rect 49193 597 49239 643
rect 49317 597 49363 643
rect 49441 597 49487 643
rect 49565 597 49611 643
rect 49689 597 49735 643
rect 49813 597 49859 643
rect 49937 597 49983 643
rect 50061 597 50107 643
rect 50185 597 50231 643
rect 50309 597 50355 643
rect 50433 597 50479 643
rect 50557 597 50603 643
rect 50681 597 50727 643
rect 50805 597 50851 643
rect 50929 597 50975 643
rect 51053 597 51099 643
rect 51177 597 51223 643
rect 51301 597 51347 643
rect 51425 597 51471 643
rect 51549 597 51595 643
rect 51673 597 51719 643
rect 51797 597 51843 643
rect 51921 597 51967 643
rect 52045 597 52091 643
rect 52169 597 52215 643
rect 52293 597 52339 643
rect 52417 597 52463 643
rect 52541 597 52587 643
rect 52665 597 52711 643
rect 52789 597 52835 643
rect 52913 597 52959 643
rect 53037 597 53083 643
rect 53161 597 53207 643
rect 53285 597 53331 643
rect 53409 597 53455 643
rect 53533 597 53579 643
rect 53657 597 53703 643
rect 53781 597 53827 643
rect 53905 597 53951 643
rect 54029 597 54075 643
rect 54153 597 54199 643
rect 54277 597 54323 643
rect 54401 597 54447 643
rect 54525 597 54571 643
rect 54649 597 54695 643
rect 54773 597 54819 643
rect 54897 597 54943 643
rect 55021 597 55067 643
rect 55145 597 55191 643
rect 55269 597 55315 643
rect 55393 597 55439 643
rect 55517 597 55563 643
rect 55641 597 55687 643
rect 55765 597 55811 643
rect 55889 597 55935 643
rect 56013 597 56059 643
rect 56137 597 56183 643
rect 56261 597 56307 643
rect 56385 597 56431 643
rect 56509 597 56555 643
rect 56633 597 56679 643
rect 56757 597 56803 643
rect 56881 597 56927 643
rect 57005 597 57051 643
rect 57129 597 57175 643
rect 57253 597 57299 643
rect 57377 597 57423 643
rect 57501 597 57547 643
rect 57625 597 57671 643
rect 57749 597 57795 643
rect 57873 597 57919 643
rect 57997 597 58043 643
rect 58121 597 58167 643
rect 58245 597 58291 643
rect 58369 597 58415 643
rect 58493 597 58539 643
rect 58617 597 58663 643
rect 58741 597 58787 643
rect 58865 597 58911 643
rect 58989 597 59035 643
rect 59113 597 59159 643
rect 59237 597 59283 643
rect 59361 597 59407 643
rect 59485 597 59531 643
rect 59609 597 59655 643
rect 59733 597 59779 643
rect 59857 597 59903 643
rect 59981 597 60027 643
rect 60105 597 60151 643
rect 60229 597 60275 643
rect 60353 597 60399 643
rect 60477 597 60523 643
rect 60601 597 60647 643
rect 60725 597 60771 643
rect 60849 597 60895 643
rect 60973 597 61019 643
rect 61097 597 61143 643
rect 61221 597 61267 643
rect 61345 597 61391 643
rect 61469 597 61515 643
rect 61593 597 61639 643
rect 61717 597 61763 643
rect 61841 597 61887 643
rect 61965 597 62011 643
rect 62089 597 62135 643
rect 62213 597 62259 643
rect 62337 597 62383 643
rect 62461 597 62507 643
rect 62585 597 62631 643
rect 62709 597 62755 643
rect 62833 597 62879 643
rect 62957 597 63003 643
rect 63081 597 63127 643
rect 63205 597 63251 643
rect 63329 597 63375 643
rect 63453 597 63499 643
rect 63577 597 63623 643
rect 63701 597 63747 643
rect 63825 597 63871 643
rect 63949 597 63995 643
rect 64073 597 64119 643
rect 64197 597 64243 643
rect 64321 597 64367 643
rect 64445 597 64491 643
rect 64569 597 64615 643
rect 64693 597 64739 643
rect 64817 597 64863 643
rect 64941 597 64987 643
rect 65065 597 65111 643
rect 65189 597 65235 643
rect 65313 597 65359 643
rect 65437 597 65483 643
rect 65561 597 65607 643
rect 65685 597 65731 643
rect 65809 597 65855 643
rect 65933 597 65979 643
rect 66057 597 66103 643
rect 66181 597 66227 643
rect 66305 597 66351 643
rect 66429 597 66475 643
rect 66553 597 66599 643
rect 66677 597 66723 643
rect 66801 597 66847 643
rect 66925 597 66971 643
rect 67049 597 67095 643
rect 67173 597 67219 643
rect 67297 597 67343 643
rect 67421 597 67467 643
rect 67545 597 67591 643
rect 67669 597 67715 643
rect 67793 597 67839 643
rect 67917 597 67963 643
rect 68041 597 68087 643
rect 68165 597 68211 643
rect 68289 597 68335 643
rect 68413 597 68459 643
rect 68537 597 68583 643
rect 68661 597 68707 643
rect 68785 597 68831 643
rect 68909 597 68955 643
rect 69033 597 69079 643
rect 69157 597 69203 643
rect 69281 597 69327 643
rect 69405 597 69451 643
rect 69529 597 69575 643
rect 69653 597 69699 643
rect 69777 597 69823 643
rect 69901 597 69947 643
rect 70025 597 70071 643
rect 70149 597 70195 643
rect 70273 597 70319 643
rect 70397 597 70443 643
rect 70521 597 70567 643
rect 70645 597 70691 643
rect 70769 597 70815 643
rect 70893 597 70939 643
rect 71017 597 71063 643
rect 71141 597 71187 643
rect 71265 597 71311 643
rect 71389 597 71435 643
rect 71513 597 71559 643
rect 71637 597 71683 643
rect 71761 597 71807 643
rect 71885 597 71931 643
rect 72009 597 72055 643
rect 72133 597 72179 643
rect 72257 597 72303 643
rect 72381 597 72427 643
rect 72505 597 72551 643
rect 72629 597 72675 643
rect 72753 597 72799 643
rect 72877 597 72923 643
rect 73001 597 73047 643
rect 73125 597 73171 643
rect 73249 597 73295 643
rect 73373 597 73419 643
rect 73497 597 73543 643
rect 73621 597 73667 643
rect 73745 597 73791 643
rect 73869 597 73915 643
rect 73993 597 74039 643
rect 74117 597 74163 643
rect 74241 597 74287 643
rect 74365 597 74411 643
rect 74489 597 74535 643
rect 74613 597 74659 643
rect 74737 597 74783 643
rect 74861 597 74907 643
rect 74985 597 75031 643
rect 75109 597 75155 643
rect 75233 597 75279 643
rect 75357 597 75403 643
rect 75481 597 75527 643
rect 75605 597 75651 643
rect 75729 597 75775 643
rect 75853 597 75899 643
rect 75977 597 76023 643
rect 76101 597 76147 643
rect 76225 597 76271 643
rect 76349 597 76395 643
rect 76473 597 76519 643
rect 76597 597 76643 643
rect 76721 597 76767 643
rect 76845 597 76891 643
rect 76969 597 77015 643
rect 77093 597 77139 643
rect 77217 597 77263 643
rect 77341 597 77387 643
rect 77465 597 77511 643
rect 77589 597 77635 643
rect 77713 597 77759 643
rect 77837 597 77883 643
rect 77961 597 78007 643
rect 78085 597 78131 643
rect 78209 597 78255 643
rect 78333 597 78379 643
rect 78457 597 78503 643
rect 78581 597 78627 643
rect 78705 597 78751 643
rect 78829 597 78875 643
rect 78953 597 78999 643
rect 79077 597 79123 643
rect 79201 597 79247 643
rect 79325 597 79371 643
rect 79449 597 79495 643
rect 79573 597 79619 643
rect 79697 597 79743 643
rect 79821 597 79867 643
rect 79945 597 79991 643
rect 80069 597 80115 643
rect 80193 597 80239 643
rect 80317 597 80363 643
rect 80441 597 80487 643
rect 80565 597 80611 643
rect 80689 597 80735 643
rect 80813 597 80859 643
rect 80937 597 80983 643
rect 81061 597 81107 643
rect 81185 597 81231 643
rect 81309 597 81355 643
rect 81433 597 81479 643
rect 81557 597 81603 643
rect 81681 597 81727 643
rect 81805 597 81851 643
rect 81929 597 81975 643
rect 82053 597 82099 643
rect 82177 597 82223 643
rect 82301 597 82347 643
rect 82425 597 82471 643
rect 82549 597 82595 643
rect 82673 597 82719 643
rect 82797 597 82843 643
rect 82921 597 82967 643
rect 83045 597 83091 643
rect 83169 597 83215 643
rect 83293 597 83339 643
rect 83417 597 83463 643
rect 83541 597 83587 643
rect 83665 597 83711 643
rect 83789 597 83835 643
rect 83913 597 83959 643
rect 84037 597 84083 643
rect 84161 597 84207 643
rect 84285 597 84331 643
rect 84409 597 84455 643
rect 84533 597 84579 643
rect 84657 597 84703 643
rect 84781 597 84827 643
rect 84905 597 84951 643
rect 85029 597 85075 643
rect 85153 597 85199 643
rect 85277 597 85323 643
rect 85401 597 85447 643
rect 85525 597 85571 643
rect 85649 597 85695 643
<< metal1 >>
rect 0 96683 85706 96694
rect 0 96637 89 96683
rect 135 96637 213 96683
rect 259 96637 337 96683
rect 383 96637 461 96683
rect 507 96637 585 96683
rect 631 96637 709 96683
rect 755 96637 833 96683
rect 879 96637 957 96683
rect 1003 96637 1081 96683
rect 1127 96637 1205 96683
rect 1251 96637 1329 96683
rect 1375 96637 1453 96683
rect 1499 96637 1577 96683
rect 1623 96637 1701 96683
rect 1747 96637 1825 96683
rect 1871 96637 1949 96683
rect 1995 96637 2073 96683
rect 2119 96637 2197 96683
rect 2243 96637 2321 96683
rect 2367 96637 2445 96683
rect 2491 96637 2569 96683
rect 2615 96637 2693 96683
rect 2739 96637 2817 96683
rect 2863 96637 2941 96683
rect 2987 96637 3065 96683
rect 3111 96637 3189 96683
rect 3235 96637 3313 96683
rect 3359 96637 3437 96683
rect 3483 96637 3561 96683
rect 3607 96637 3685 96683
rect 3731 96637 3809 96683
rect 3855 96637 3933 96683
rect 3979 96637 4057 96683
rect 4103 96637 4181 96683
rect 4227 96637 4305 96683
rect 4351 96637 4429 96683
rect 4475 96637 4553 96683
rect 4599 96637 4677 96683
rect 4723 96637 4801 96683
rect 4847 96637 4925 96683
rect 4971 96637 5049 96683
rect 5095 96637 5173 96683
rect 5219 96637 5297 96683
rect 5343 96637 5421 96683
rect 5467 96637 5545 96683
rect 5591 96637 5669 96683
rect 5715 96637 5793 96683
rect 5839 96637 5917 96683
rect 5963 96637 6041 96683
rect 6087 96637 6165 96683
rect 6211 96637 6289 96683
rect 6335 96637 6413 96683
rect 6459 96637 6537 96683
rect 6583 96637 6661 96683
rect 6707 96637 6785 96683
rect 6831 96637 6909 96683
rect 6955 96637 7033 96683
rect 7079 96637 7157 96683
rect 7203 96637 7281 96683
rect 7327 96637 7405 96683
rect 7451 96637 7529 96683
rect 7575 96637 7653 96683
rect 7699 96637 7777 96683
rect 7823 96637 7901 96683
rect 7947 96637 8025 96683
rect 8071 96637 8149 96683
rect 8195 96637 8273 96683
rect 8319 96637 8397 96683
rect 8443 96637 8521 96683
rect 8567 96637 8645 96683
rect 8691 96637 8769 96683
rect 8815 96637 8893 96683
rect 8939 96637 9017 96683
rect 9063 96637 9141 96683
rect 9187 96637 9265 96683
rect 9311 96637 9389 96683
rect 9435 96637 9513 96683
rect 9559 96637 9637 96683
rect 9683 96637 9761 96683
rect 9807 96637 9885 96683
rect 9931 96637 10009 96683
rect 10055 96637 10133 96683
rect 10179 96637 10257 96683
rect 10303 96637 10381 96683
rect 10427 96637 10505 96683
rect 10551 96637 10629 96683
rect 10675 96637 10753 96683
rect 10799 96637 10877 96683
rect 10923 96637 11001 96683
rect 11047 96637 11125 96683
rect 11171 96637 11249 96683
rect 11295 96637 11373 96683
rect 11419 96637 11497 96683
rect 11543 96637 11621 96683
rect 11667 96637 11745 96683
rect 11791 96637 11869 96683
rect 11915 96637 11993 96683
rect 12039 96637 12117 96683
rect 12163 96637 12241 96683
rect 12287 96637 12365 96683
rect 12411 96637 12489 96683
rect 12535 96637 12613 96683
rect 12659 96637 12737 96683
rect 12783 96637 12861 96683
rect 12907 96637 12985 96683
rect 13031 96637 13109 96683
rect 13155 96637 13233 96683
rect 13279 96637 13357 96683
rect 13403 96637 13481 96683
rect 13527 96637 13605 96683
rect 13651 96637 13729 96683
rect 13775 96637 13853 96683
rect 13899 96637 13977 96683
rect 14023 96637 14101 96683
rect 14147 96637 14225 96683
rect 14271 96637 14349 96683
rect 14395 96637 14473 96683
rect 14519 96637 14597 96683
rect 14643 96637 14721 96683
rect 14767 96637 14845 96683
rect 14891 96637 14969 96683
rect 15015 96637 15093 96683
rect 15139 96637 15217 96683
rect 15263 96637 15341 96683
rect 15387 96637 15465 96683
rect 15511 96637 15589 96683
rect 15635 96637 15713 96683
rect 15759 96637 15837 96683
rect 15883 96637 15961 96683
rect 16007 96637 16085 96683
rect 16131 96637 16209 96683
rect 16255 96637 16333 96683
rect 16379 96637 16457 96683
rect 16503 96637 16581 96683
rect 16627 96637 16705 96683
rect 16751 96637 16829 96683
rect 16875 96637 16953 96683
rect 16999 96637 17077 96683
rect 17123 96637 17201 96683
rect 17247 96637 17325 96683
rect 17371 96637 17449 96683
rect 17495 96637 17573 96683
rect 17619 96637 17697 96683
rect 17743 96637 17821 96683
rect 17867 96637 17945 96683
rect 17991 96637 18069 96683
rect 18115 96637 18193 96683
rect 18239 96637 18317 96683
rect 18363 96637 18441 96683
rect 18487 96637 18565 96683
rect 18611 96637 18689 96683
rect 18735 96637 18813 96683
rect 18859 96637 18937 96683
rect 18983 96637 19061 96683
rect 19107 96637 19185 96683
rect 19231 96637 19309 96683
rect 19355 96637 19433 96683
rect 19479 96637 19557 96683
rect 19603 96637 19681 96683
rect 19727 96637 19805 96683
rect 19851 96637 19929 96683
rect 19975 96637 20053 96683
rect 20099 96637 20177 96683
rect 20223 96637 20301 96683
rect 20347 96637 20425 96683
rect 20471 96637 20549 96683
rect 20595 96637 20673 96683
rect 20719 96637 20797 96683
rect 20843 96637 20921 96683
rect 20967 96637 21045 96683
rect 21091 96637 21169 96683
rect 21215 96637 21293 96683
rect 21339 96637 21417 96683
rect 21463 96637 21541 96683
rect 21587 96637 21665 96683
rect 21711 96637 21789 96683
rect 21835 96637 21913 96683
rect 21959 96637 22037 96683
rect 22083 96637 22161 96683
rect 22207 96637 22285 96683
rect 22331 96637 22409 96683
rect 22455 96637 22533 96683
rect 22579 96637 22657 96683
rect 22703 96637 22781 96683
rect 22827 96637 22905 96683
rect 22951 96637 23029 96683
rect 23075 96637 23153 96683
rect 23199 96637 23277 96683
rect 23323 96637 23401 96683
rect 23447 96637 23525 96683
rect 23571 96637 23649 96683
rect 23695 96637 23773 96683
rect 23819 96637 23897 96683
rect 23943 96637 24021 96683
rect 24067 96637 24145 96683
rect 24191 96637 24269 96683
rect 24315 96637 24393 96683
rect 24439 96637 24517 96683
rect 24563 96637 24641 96683
rect 24687 96637 24765 96683
rect 24811 96637 24889 96683
rect 24935 96637 25013 96683
rect 25059 96637 25137 96683
rect 25183 96637 25261 96683
rect 25307 96637 25385 96683
rect 25431 96637 25509 96683
rect 25555 96637 25633 96683
rect 25679 96637 25757 96683
rect 25803 96637 25881 96683
rect 25927 96637 26005 96683
rect 26051 96637 26129 96683
rect 26175 96637 26253 96683
rect 26299 96637 26377 96683
rect 26423 96637 26501 96683
rect 26547 96637 26625 96683
rect 26671 96637 26749 96683
rect 26795 96637 26873 96683
rect 26919 96637 26997 96683
rect 27043 96637 27121 96683
rect 27167 96637 27245 96683
rect 27291 96637 27369 96683
rect 27415 96637 27493 96683
rect 27539 96637 27617 96683
rect 27663 96637 27741 96683
rect 27787 96637 27865 96683
rect 27911 96637 27989 96683
rect 28035 96637 28113 96683
rect 28159 96637 28237 96683
rect 28283 96637 28361 96683
rect 28407 96637 28485 96683
rect 28531 96637 28609 96683
rect 28655 96637 28733 96683
rect 28779 96637 28857 96683
rect 28903 96637 28981 96683
rect 29027 96637 29105 96683
rect 29151 96637 29229 96683
rect 29275 96637 29353 96683
rect 29399 96637 29477 96683
rect 29523 96637 29601 96683
rect 29647 96637 29725 96683
rect 29771 96637 29849 96683
rect 29895 96637 29973 96683
rect 30019 96637 30097 96683
rect 30143 96637 30221 96683
rect 30267 96637 30345 96683
rect 30391 96637 30469 96683
rect 30515 96637 30593 96683
rect 30639 96637 30717 96683
rect 30763 96637 30841 96683
rect 30887 96637 30965 96683
rect 31011 96637 31089 96683
rect 31135 96637 31213 96683
rect 31259 96637 31337 96683
rect 31383 96637 31461 96683
rect 31507 96637 31585 96683
rect 31631 96637 31709 96683
rect 31755 96637 31833 96683
rect 31879 96637 31957 96683
rect 32003 96637 32081 96683
rect 32127 96637 32205 96683
rect 32251 96637 32329 96683
rect 32375 96637 32453 96683
rect 32499 96637 32577 96683
rect 32623 96637 32701 96683
rect 32747 96637 32825 96683
rect 32871 96637 32949 96683
rect 32995 96637 33073 96683
rect 33119 96637 33197 96683
rect 33243 96637 33321 96683
rect 33367 96637 33445 96683
rect 33491 96637 33569 96683
rect 33615 96637 33693 96683
rect 33739 96637 33817 96683
rect 33863 96637 33941 96683
rect 33987 96637 34065 96683
rect 34111 96637 34189 96683
rect 34235 96637 34313 96683
rect 34359 96637 34437 96683
rect 34483 96637 34561 96683
rect 34607 96637 34685 96683
rect 34731 96637 34809 96683
rect 34855 96637 34933 96683
rect 34979 96637 35057 96683
rect 35103 96637 35181 96683
rect 35227 96637 35305 96683
rect 35351 96637 35429 96683
rect 35475 96637 35553 96683
rect 35599 96637 35677 96683
rect 35723 96637 35801 96683
rect 35847 96637 35925 96683
rect 35971 96637 36049 96683
rect 36095 96637 36173 96683
rect 36219 96637 36297 96683
rect 36343 96637 36421 96683
rect 36467 96637 36545 96683
rect 36591 96637 36669 96683
rect 36715 96637 36793 96683
rect 36839 96637 36917 96683
rect 36963 96637 37041 96683
rect 37087 96637 37165 96683
rect 37211 96637 37289 96683
rect 37335 96637 37413 96683
rect 37459 96637 37537 96683
rect 37583 96637 37661 96683
rect 37707 96637 37785 96683
rect 37831 96637 37909 96683
rect 37955 96637 38033 96683
rect 38079 96637 38157 96683
rect 38203 96637 38281 96683
rect 38327 96637 38405 96683
rect 38451 96637 38529 96683
rect 38575 96637 38653 96683
rect 38699 96637 38777 96683
rect 38823 96637 38901 96683
rect 38947 96637 39025 96683
rect 39071 96637 39149 96683
rect 39195 96637 39273 96683
rect 39319 96637 39397 96683
rect 39443 96637 39521 96683
rect 39567 96637 39645 96683
rect 39691 96637 39769 96683
rect 39815 96637 39893 96683
rect 39939 96637 40017 96683
rect 40063 96637 40141 96683
rect 40187 96637 40265 96683
rect 40311 96637 40389 96683
rect 40435 96637 40513 96683
rect 40559 96637 40637 96683
rect 40683 96637 40761 96683
rect 40807 96637 40885 96683
rect 40931 96637 41009 96683
rect 41055 96637 41133 96683
rect 41179 96637 41257 96683
rect 41303 96637 41381 96683
rect 41427 96637 41505 96683
rect 41551 96637 41629 96683
rect 41675 96637 41753 96683
rect 41799 96637 41877 96683
rect 41923 96637 42001 96683
rect 42047 96637 42125 96683
rect 42171 96637 42249 96683
rect 42295 96637 42373 96683
rect 42419 96637 42497 96683
rect 42543 96637 42621 96683
rect 42667 96637 42745 96683
rect 42791 96637 42869 96683
rect 42915 96637 42993 96683
rect 43039 96637 43117 96683
rect 43163 96637 43241 96683
rect 43287 96637 43365 96683
rect 43411 96637 43489 96683
rect 43535 96637 43613 96683
rect 43659 96637 43737 96683
rect 43783 96637 43861 96683
rect 43907 96637 43985 96683
rect 44031 96637 44109 96683
rect 44155 96637 44233 96683
rect 44279 96637 44357 96683
rect 44403 96637 44481 96683
rect 44527 96637 44605 96683
rect 44651 96637 44729 96683
rect 44775 96637 44853 96683
rect 44899 96637 44977 96683
rect 45023 96637 45101 96683
rect 45147 96637 45225 96683
rect 45271 96637 45349 96683
rect 45395 96637 45473 96683
rect 45519 96637 45597 96683
rect 45643 96637 45721 96683
rect 45767 96637 45845 96683
rect 45891 96637 45969 96683
rect 46015 96637 46093 96683
rect 46139 96637 46217 96683
rect 46263 96637 46341 96683
rect 46387 96637 46465 96683
rect 46511 96637 46589 96683
rect 46635 96637 46713 96683
rect 46759 96637 46837 96683
rect 46883 96637 46961 96683
rect 47007 96637 47085 96683
rect 47131 96637 47209 96683
rect 47255 96637 47333 96683
rect 47379 96637 47457 96683
rect 47503 96637 47581 96683
rect 47627 96637 47705 96683
rect 47751 96637 47829 96683
rect 47875 96637 47953 96683
rect 47999 96637 48077 96683
rect 48123 96637 48201 96683
rect 48247 96637 48325 96683
rect 48371 96637 48449 96683
rect 48495 96637 48573 96683
rect 48619 96637 48697 96683
rect 48743 96637 48821 96683
rect 48867 96637 48945 96683
rect 48991 96637 49069 96683
rect 49115 96637 49193 96683
rect 49239 96637 49317 96683
rect 49363 96637 49441 96683
rect 49487 96637 49565 96683
rect 49611 96637 49689 96683
rect 49735 96637 49813 96683
rect 49859 96637 49937 96683
rect 49983 96637 50061 96683
rect 50107 96637 50185 96683
rect 50231 96637 50309 96683
rect 50355 96637 50433 96683
rect 50479 96637 50557 96683
rect 50603 96637 50681 96683
rect 50727 96637 50805 96683
rect 50851 96637 50929 96683
rect 50975 96637 51053 96683
rect 51099 96637 51177 96683
rect 51223 96637 51301 96683
rect 51347 96637 51425 96683
rect 51471 96637 51549 96683
rect 51595 96637 51673 96683
rect 51719 96637 51797 96683
rect 51843 96637 51921 96683
rect 51967 96637 52045 96683
rect 52091 96637 52169 96683
rect 52215 96637 52293 96683
rect 52339 96637 52417 96683
rect 52463 96637 52541 96683
rect 52587 96637 52665 96683
rect 52711 96637 52789 96683
rect 52835 96637 52913 96683
rect 52959 96637 53037 96683
rect 53083 96637 53161 96683
rect 53207 96637 53285 96683
rect 53331 96637 53409 96683
rect 53455 96637 53533 96683
rect 53579 96637 53657 96683
rect 53703 96637 53781 96683
rect 53827 96637 53905 96683
rect 53951 96637 54029 96683
rect 54075 96637 54153 96683
rect 54199 96637 54277 96683
rect 54323 96637 54401 96683
rect 54447 96637 54525 96683
rect 54571 96637 54649 96683
rect 54695 96637 54773 96683
rect 54819 96637 54897 96683
rect 54943 96637 55021 96683
rect 55067 96637 55145 96683
rect 55191 96637 55269 96683
rect 55315 96637 55393 96683
rect 55439 96637 55517 96683
rect 55563 96637 55641 96683
rect 55687 96637 55765 96683
rect 55811 96637 55889 96683
rect 55935 96637 56013 96683
rect 56059 96637 56137 96683
rect 56183 96637 56261 96683
rect 56307 96637 56385 96683
rect 56431 96637 56509 96683
rect 56555 96637 56633 96683
rect 56679 96637 56757 96683
rect 56803 96637 56881 96683
rect 56927 96637 57005 96683
rect 57051 96637 57129 96683
rect 57175 96637 57253 96683
rect 57299 96637 57377 96683
rect 57423 96637 57501 96683
rect 57547 96637 57625 96683
rect 57671 96637 57749 96683
rect 57795 96637 57873 96683
rect 57919 96637 57997 96683
rect 58043 96637 58121 96683
rect 58167 96637 58245 96683
rect 58291 96637 58369 96683
rect 58415 96637 58493 96683
rect 58539 96637 58617 96683
rect 58663 96637 58741 96683
rect 58787 96637 58865 96683
rect 58911 96637 58989 96683
rect 59035 96637 59113 96683
rect 59159 96637 59237 96683
rect 59283 96637 59361 96683
rect 59407 96637 59485 96683
rect 59531 96637 59609 96683
rect 59655 96637 59733 96683
rect 59779 96637 59857 96683
rect 59903 96637 59981 96683
rect 60027 96637 60105 96683
rect 60151 96637 60229 96683
rect 60275 96637 60353 96683
rect 60399 96637 60477 96683
rect 60523 96637 60601 96683
rect 60647 96637 60725 96683
rect 60771 96637 60849 96683
rect 60895 96637 60973 96683
rect 61019 96637 61097 96683
rect 61143 96637 61221 96683
rect 61267 96637 61345 96683
rect 61391 96637 61469 96683
rect 61515 96637 61593 96683
rect 61639 96637 61717 96683
rect 61763 96637 61841 96683
rect 61887 96637 61965 96683
rect 62011 96637 62089 96683
rect 62135 96637 62213 96683
rect 62259 96637 62337 96683
rect 62383 96637 62461 96683
rect 62507 96637 62585 96683
rect 62631 96637 62709 96683
rect 62755 96637 62833 96683
rect 62879 96637 62957 96683
rect 63003 96637 63081 96683
rect 63127 96637 63205 96683
rect 63251 96637 63329 96683
rect 63375 96637 63453 96683
rect 63499 96637 63577 96683
rect 63623 96637 63701 96683
rect 63747 96637 63825 96683
rect 63871 96637 63949 96683
rect 63995 96637 64073 96683
rect 64119 96637 64197 96683
rect 64243 96637 64321 96683
rect 64367 96637 64445 96683
rect 64491 96637 64569 96683
rect 64615 96637 64693 96683
rect 64739 96637 64817 96683
rect 64863 96637 64941 96683
rect 64987 96637 65065 96683
rect 65111 96637 65189 96683
rect 65235 96637 65313 96683
rect 65359 96637 65437 96683
rect 65483 96637 65561 96683
rect 65607 96637 65685 96683
rect 65731 96637 65809 96683
rect 65855 96637 65933 96683
rect 65979 96637 66057 96683
rect 66103 96637 66181 96683
rect 66227 96637 66305 96683
rect 66351 96637 66429 96683
rect 66475 96637 66553 96683
rect 66599 96637 66677 96683
rect 66723 96637 66801 96683
rect 66847 96637 66925 96683
rect 66971 96637 67049 96683
rect 67095 96637 67173 96683
rect 67219 96637 67297 96683
rect 67343 96637 67421 96683
rect 67467 96637 67545 96683
rect 67591 96637 67669 96683
rect 67715 96637 67793 96683
rect 67839 96637 67917 96683
rect 67963 96637 68041 96683
rect 68087 96637 68165 96683
rect 68211 96637 68289 96683
rect 68335 96637 68413 96683
rect 68459 96637 68537 96683
rect 68583 96637 68661 96683
rect 68707 96637 68785 96683
rect 68831 96637 68909 96683
rect 68955 96637 69033 96683
rect 69079 96637 69157 96683
rect 69203 96637 69281 96683
rect 69327 96637 69405 96683
rect 69451 96637 69529 96683
rect 69575 96637 69653 96683
rect 69699 96637 69777 96683
rect 69823 96637 69901 96683
rect 69947 96637 70025 96683
rect 70071 96637 70149 96683
rect 70195 96637 70273 96683
rect 70319 96637 70397 96683
rect 70443 96637 70521 96683
rect 70567 96637 70645 96683
rect 70691 96637 70769 96683
rect 70815 96637 70893 96683
rect 70939 96637 71017 96683
rect 71063 96637 71141 96683
rect 71187 96637 71265 96683
rect 71311 96637 71389 96683
rect 71435 96637 71513 96683
rect 71559 96637 71637 96683
rect 71683 96637 71761 96683
rect 71807 96637 71885 96683
rect 71931 96637 72009 96683
rect 72055 96637 72133 96683
rect 72179 96637 72257 96683
rect 72303 96637 72381 96683
rect 72427 96637 72505 96683
rect 72551 96637 72629 96683
rect 72675 96637 72753 96683
rect 72799 96637 72877 96683
rect 72923 96637 73001 96683
rect 73047 96637 73125 96683
rect 73171 96637 73249 96683
rect 73295 96637 73373 96683
rect 73419 96637 73497 96683
rect 73543 96637 73621 96683
rect 73667 96637 73745 96683
rect 73791 96637 73869 96683
rect 73915 96637 73993 96683
rect 74039 96637 74117 96683
rect 74163 96637 74241 96683
rect 74287 96637 74365 96683
rect 74411 96637 74489 96683
rect 74535 96637 74613 96683
rect 74659 96637 74737 96683
rect 74783 96637 74861 96683
rect 74907 96637 74985 96683
rect 75031 96637 75109 96683
rect 75155 96637 75233 96683
rect 75279 96637 75357 96683
rect 75403 96637 75481 96683
rect 75527 96637 75605 96683
rect 75651 96637 75729 96683
rect 75775 96637 75853 96683
rect 75899 96637 75977 96683
rect 76023 96637 76101 96683
rect 76147 96637 76225 96683
rect 76271 96637 76349 96683
rect 76395 96637 76473 96683
rect 76519 96637 76597 96683
rect 76643 96637 76721 96683
rect 76767 96637 76845 96683
rect 76891 96637 76969 96683
rect 77015 96637 77093 96683
rect 77139 96637 77217 96683
rect 77263 96637 77341 96683
rect 77387 96637 77465 96683
rect 77511 96637 77589 96683
rect 77635 96637 77713 96683
rect 77759 96637 77837 96683
rect 77883 96637 77961 96683
rect 78007 96637 78085 96683
rect 78131 96637 78209 96683
rect 78255 96637 78333 96683
rect 78379 96637 78457 96683
rect 78503 96637 78581 96683
rect 78627 96637 78705 96683
rect 78751 96637 78829 96683
rect 78875 96637 78953 96683
rect 78999 96637 79077 96683
rect 79123 96637 79201 96683
rect 79247 96637 79325 96683
rect 79371 96637 79449 96683
rect 79495 96637 79573 96683
rect 79619 96637 79697 96683
rect 79743 96637 79821 96683
rect 79867 96637 79945 96683
rect 79991 96637 80069 96683
rect 80115 96637 80193 96683
rect 80239 96637 80317 96683
rect 80363 96637 80441 96683
rect 80487 96637 80565 96683
rect 80611 96637 80689 96683
rect 80735 96637 80813 96683
rect 80859 96637 80937 96683
rect 80983 96637 81061 96683
rect 81107 96637 81185 96683
rect 81231 96637 81309 96683
rect 81355 96637 81433 96683
rect 81479 96637 81557 96683
rect 81603 96637 81681 96683
rect 81727 96637 81805 96683
rect 81851 96637 81929 96683
rect 81975 96637 82053 96683
rect 82099 96637 82177 96683
rect 82223 96637 82301 96683
rect 82347 96637 82425 96683
rect 82471 96637 82549 96683
rect 82595 96637 82673 96683
rect 82719 96637 82797 96683
rect 82843 96637 82921 96683
rect 82967 96637 83045 96683
rect 83091 96637 83169 96683
rect 83215 96637 83293 96683
rect 83339 96637 83417 96683
rect 83463 96637 83541 96683
rect 83587 96637 83665 96683
rect 83711 96637 83789 96683
rect 83835 96637 83913 96683
rect 83959 96637 84037 96683
rect 84083 96637 84161 96683
rect 84207 96637 84285 96683
rect 84331 96637 84409 96683
rect 84455 96637 84533 96683
rect 84579 96637 84657 96683
rect 84703 96637 84781 96683
rect 84827 96637 84905 96683
rect 84951 96637 85029 96683
rect 85075 96637 85153 96683
rect 85199 96637 85277 96683
rect 85323 96637 85401 96683
rect 85447 96637 85525 96683
rect 85571 96637 85649 96683
rect 85695 96637 85706 96683
rect 0 96559 85706 96637
rect 0 96513 89 96559
rect 135 96513 213 96559
rect 259 96513 337 96559
rect 383 96513 461 96559
rect 507 96513 585 96559
rect 631 96513 709 96559
rect 755 96513 833 96559
rect 879 96513 957 96559
rect 1003 96513 1081 96559
rect 1127 96513 1205 96559
rect 1251 96513 1329 96559
rect 1375 96513 1453 96559
rect 1499 96513 1577 96559
rect 1623 96513 1701 96559
rect 1747 96513 1825 96559
rect 1871 96513 1949 96559
rect 1995 96513 2073 96559
rect 2119 96513 2197 96559
rect 2243 96513 2321 96559
rect 2367 96513 2445 96559
rect 2491 96513 2569 96559
rect 2615 96513 2693 96559
rect 2739 96513 2817 96559
rect 2863 96513 2941 96559
rect 2987 96513 3065 96559
rect 3111 96513 3189 96559
rect 3235 96513 3313 96559
rect 3359 96513 3437 96559
rect 3483 96513 3561 96559
rect 3607 96513 3685 96559
rect 3731 96513 3809 96559
rect 3855 96513 3933 96559
rect 3979 96513 4057 96559
rect 4103 96513 4181 96559
rect 4227 96513 4305 96559
rect 4351 96513 4429 96559
rect 4475 96513 4553 96559
rect 4599 96513 4677 96559
rect 4723 96513 4801 96559
rect 4847 96513 4925 96559
rect 4971 96513 5049 96559
rect 5095 96513 5173 96559
rect 5219 96513 5297 96559
rect 5343 96513 5421 96559
rect 5467 96513 5545 96559
rect 5591 96513 5669 96559
rect 5715 96513 5793 96559
rect 5839 96513 5917 96559
rect 5963 96513 6041 96559
rect 6087 96513 6165 96559
rect 6211 96513 6289 96559
rect 6335 96513 6413 96559
rect 6459 96513 6537 96559
rect 6583 96513 6661 96559
rect 6707 96513 6785 96559
rect 6831 96513 6909 96559
rect 6955 96513 7033 96559
rect 7079 96513 7157 96559
rect 7203 96513 7281 96559
rect 7327 96513 7405 96559
rect 7451 96513 7529 96559
rect 7575 96513 7653 96559
rect 7699 96513 7777 96559
rect 7823 96513 7901 96559
rect 7947 96513 8025 96559
rect 8071 96513 8149 96559
rect 8195 96513 8273 96559
rect 8319 96513 8397 96559
rect 8443 96513 8521 96559
rect 8567 96513 8645 96559
rect 8691 96513 8769 96559
rect 8815 96513 8893 96559
rect 8939 96513 9017 96559
rect 9063 96513 9141 96559
rect 9187 96513 9265 96559
rect 9311 96513 9389 96559
rect 9435 96513 9513 96559
rect 9559 96513 9637 96559
rect 9683 96513 9761 96559
rect 9807 96513 9885 96559
rect 9931 96513 10009 96559
rect 10055 96513 10133 96559
rect 10179 96513 10257 96559
rect 10303 96513 10381 96559
rect 10427 96513 10505 96559
rect 10551 96513 10629 96559
rect 10675 96513 10753 96559
rect 10799 96513 10877 96559
rect 10923 96513 11001 96559
rect 11047 96513 11125 96559
rect 11171 96513 11249 96559
rect 11295 96513 11373 96559
rect 11419 96513 11497 96559
rect 11543 96513 11621 96559
rect 11667 96513 11745 96559
rect 11791 96513 11869 96559
rect 11915 96513 11993 96559
rect 12039 96513 12117 96559
rect 12163 96513 12241 96559
rect 12287 96513 12365 96559
rect 12411 96513 12489 96559
rect 12535 96513 12613 96559
rect 12659 96513 12737 96559
rect 12783 96513 12861 96559
rect 12907 96513 12985 96559
rect 13031 96513 13109 96559
rect 13155 96513 13233 96559
rect 13279 96513 13357 96559
rect 13403 96513 13481 96559
rect 13527 96513 13605 96559
rect 13651 96513 13729 96559
rect 13775 96513 13853 96559
rect 13899 96513 13977 96559
rect 14023 96513 14101 96559
rect 14147 96513 14225 96559
rect 14271 96513 14349 96559
rect 14395 96513 14473 96559
rect 14519 96513 14597 96559
rect 14643 96513 14721 96559
rect 14767 96513 14845 96559
rect 14891 96513 14969 96559
rect 15015 96513 15093 96559
rect 15139 96513 15217 96559
rect 15263 96513 15341 96559
rect 15387 96513 15465 96559
rect 15511 96513 15589 96559
rect 15635 96513 15713 96559
rect 15759 96513 15837 96559
rect 15883 96513 15961 96559
rect 16007 96513 16085 96559
rect 16131 96513 16209 96559
rect 16255 96513 16333 96559
rect 16379 96513 16457 96559
rect 16503 96513 16581 96559
rect 16627 96513 16705 96559
rect 16751 96513 16829 96559
rect 16875 96513 16953 96559
rect 16999 96513 17077 96559
rect 17123 96513 17201 96559
rect 17247 96513 17325 96559
rect 17371 96513 17449 96559
rect 17495 96513 17573 96559
rect 17619 96513 17697 96559
rect 17743 96513 17821 96559
rect 17867 96513 17945 96559
rect 17991 96513 18069 96559
rect 18115 96513 18193 96559
rect 18239 96513 18317 96559
rect 18363 96513 18441 96559
rect 18487 96513 18565 96559
rect 18611 96513 18689 96559
rect 18735 96513 18813 96559
rect 18859 96513 18937 96559
rect 18983 96513 19061 96559
rect 19107 96513 19185 96559
rect 19231 96513 19309 96559
rect 19355 96513 19433 96559
rect 19479 96513 19557 96559
rect 19603 96513 19681 96559
rect 19727 96513 19805 96559
rect 19851 96513 19929 96559
rect 19975 96513 20053 96559
rect 20099 96513 20177 96559
rect 20223 96513 20301 96559
rect 20347 96513 20425 96559
rect 20471 96513 20549 96559
rect 20595 96513 20673 96559
rect 20719 96513 20797 96559
rect 20843 96513 20921 96559
rect 20967 96513 21045 96559
rect 21091 96513 21169 96559
rect 21215 96513 21293 96559
rect 21339 96513 21417 96559
rect 21463 96513 21541 96559
rect 21587 96513 21665 96559
rect 21711 96513 21789 96559
rect 21835 96513 21913 96559
rect 21959 96513 22037 96559
rect 22083 96513 22161 96559
rect 22207 96513 22285 96559
rect 22331 96513 22409 96559
rect 22455 96513 22533 96559
rect 22579 96513 22657 96559
rect 22703 96513 22781 96559
rect 22827 96513 22905 96559
rect 22951 96513 23029 96559
rect 23075 96513 23153 96559
rect 23199 96513 23277 96559
rect 23323 96513 23401 96559
rect 23447 96513 23525 96559
rect 23571 96513 23649 96559
rect 23695 96513 23773 96559
rect 23819 96513 23897 96559
rect 23943 96513 24021 96559
rect 24067 96513 24145 96559
rect 24191 96513 24269 96559
rect 24315 96513 24393 96559
rect 24439 96513 24517 96559
rect 24563 96513 24641 96559
rect 24687 96513 24765 96559
rect 24811 96513 24889 96559
rect 24935 96513 25013 96559
rect 25059 96513 25137 96559
rect 25183 96513 25261 96559
rect 25307 96513 25385 96559
rect 25431 96513 25509 96559
rect 25555 96513 25633 96559
rect 25679 96513 25757 96559
rect 25803 96513 25881 96559
rect 25927 96513 26005 96559
rect 26051 96513 26129 96559
rect 26175 96513 26253 96559
rect 26299 96513 26377 96559
rect 26423 96513 26501 96559
rect 26547 96513 26625 96559
rect 26671 96513 26749 96559
rect 26795 96513 26873 96559
rect 26919 96513 26997 96559
rect 27043 96513 27121 96559
rect 27167 96513 27245 96559
rect 27291 96513 27369 96559
rect 27415 96513 27493 96559
rect 27539 96513 27617 96559
rect 27663 96513 27741 96559
rect 27787 96513 27865 96559
rect 27911 96513 27989 96559
rect 28035 96513 28113 96559
rect 28159 96513 28237 96559
rect 28283 96513 28361 96559
rect 28407 96513 28485 96559
rect 28531 96513 28609 96559
rect 28655 96513 28733 96559
rect 28779 96513 28857 96559
rect 28903 96513 28981 96559
rect 29027 96513 29105 96559
rect 29151 96513 29229 96559
rect 29275 96513 29353 96559
rect 29399 96513 29477 96559
rect 29523 96513 29601 96559
rect 29647 96513 29725 96559
rect 29771 96513 29849 96559
rect 29895 96513 29973 96559
rect 30019 96513 30097 96559
rect 30143 96513 30221 96559
rect 30267 96513 30345 96559
rect 30391 96513 30469 96559
rect 30515 96513 30593 96559
rect 30639 96513 30717 96559
rect 30763 96513 30841 96559
rect 30887 96513 30965 96559
rect 31011 96513 31089 96559
rect 31135 96513 31213 96559
rect 31259 96513 31337 96559
rect 31383 96513 31461 96559
rect 31507 96513 31585 96559
rect 31631 96513 31709 96559
rect 31755 96513 31833 96559
rect 31879 96513 31957 96559
rect 32003 96513 32081 96559
rect 32127 96513 32205 96559
rect 32251 96513 32329 96559
rect 32375 96513 32453 96559
rect 32499 96513 32577 96559
rect 32623 96513 32701 96559
rect 32747 96513 32825 96559
rect 32871 96513 32949 96559
rect 32995 96513 33073 96559
rect 33119 96513 33197 96559
rect 33243 96513 33321 96559
rect 33367 96513 33445 96559
rect 33491 96513 33569 96559
rect 33615 96513 33693 96559
rect 33739 96513 33817 96559
rect 33863 96513 33941 96559
rect 33987 96513 34065 96559
rect 34111 96513 34189 96559
rect 34235 96513 34313 96559
rect 34359 96513 34437 96559
rect 34483 96513 34561 96559
rect 34607 96513 34685 96559
rect 34731 96513 34809 96559
rect 34855 96513 34933 96559
rect 34979 96513 35057 96559
rect 35103 96513 35181 96559
rect 35227 96513 35305 96559
rect 35351 96513 35429 96559
rect 35475 96513 35553 96559
rect 35599 96513 35677 96559
rect 35723 96513 35801 96559
rect 35847 96513 35925 96559
rect 35971 96513 36049 96559
rect 36095 96513 36173 96559
rect 36219 96513 36297 96559
rect 36343 96513 36421 96559
rect 36467 96513 36545 96559
rect 36591 96513 36669 96559
rect 36715 96513 36793 96559
rect 36839 96513 36917 96559
rect 36963 96513 37041 96559
rect 37087 96513 37165 96559
rect 37211 96513 37289 96559
rect 37335 96513 37413 96559
rect 37459 96513 37537 96559
rect 37583 96513 37661 96559
rect 37707 96513 37785 96559
rect 37831 96513 37909 96559
rect 37955 96513 38033 96559
rect 38079 96513 38157 96559
rect 38203 96513 38281 96559
rect 38327 96513 38405 96559
rect 38451 96513 38529 96559
rect 38575 96513 38653 96559
rect 38699 96513 38777 96559
rect 38823 96513 38901 96559
rect 38947 96513 39025 96559
rect 39071 96513 39149 96559
rect 39195 96513 39273 96559
rect 39319 96513 39397 96559
rect 39443 96513 39521 96559
rect 39567 96513 39645 96559
rect 39691 96513 39769 96559
rect 39815 96513 39893 96559
rect 39939 96513 40017 96559
rect 40063 96513 40141 96559
rect 40187 96513 40265 96559
rect 40311 96513 40389 96559
rect 40435 96513 40513 96559
rect 40559 96513 40637 96559
rect 40683 96513 40761 96559
rect 40807 96513 40885 96559
rect 40931 96513 41009 96559
rect 41055 96513 41133 96559
rect 41179 96513 41257 96559
rect 41303 96513 41381 96559
rect 41427 96513 41505 96559
rect 41551 96513 41629 96559
rect 41675 96513 41753 96559
rect 41799 96513 41877 96559
rect 41923 96513 42001 96559
rect 42047 96513 42125 96559
rect 42171 96513 42249 96559
rect 42295 96513 42373 96559
rect 42419 96513 42497 96559
rect 42543 96513 42621 96559
rect 42667 96513 42745 96559
rect 42791 96513 42869 96559
rect 42915 96513 42993 96559
rect 43039 96513 43117 96559
rect 43163 96513 43241 96559
rect 43287 96513 43365 96559
rect 43411 96513 43489 96559
rect 43535 96513 43613 96559
rect 43659 96513 43737 96559
rect 43783 96513 43861 96559
rect 43907 96513 43985 96559
rect 44031 96513 44109 96559
rect 44155 96513 44233 96559
rect 44279 96513 44357 96559
rect 44403 96513 44481 96559
rect 44527 96513 44605 96559
rect 44651 96513 44729 96559
rect 44775 96513 44853 96559
rect 44899 96513 44977 96559
rect 45023 96513 45101 96559
rect 45147 96513 45225 96559
rect 45271 96513 45349 96559
rect 45395 96513 45473 96559
rect 45519 96513 45597 96559
rect 45643 96513 45721 96559
rect 45767 96513 45845 96559
rect 45891 96513 45969 96559
rect 46015 96513 46093 96559
rect 46139 96513 46217 96559
rect 46263 96513 46341 96559
rect 46387 96513 46465 96559
rect 46511 96513 46589 96559
rect 46635 96513 46713 96559
rect 46759 96513 46837 96559
rect 46883 96513 46961 96559
rect 47007 96513 47085 96559
rect 47131 96513 47209 96559
rect 47255 96513 47333 96559
rect 47379 96513 47457 96559
rect 47503 96513 47581 96559
rect 47627 96513 47705 96559
rect 47751 96513 47829 96559
rect 47875 96513 47953 96559
rect 47999 96513 48077 96559
rect 48123 96513 48201 96559
rect 48247 96513 48325 96559
rect 48371 96513 48449 96559
rect 48495 96513 48573 96559
rect 48619 96513 48697 96559
rect 48743 96513 48821 96559
rect 48867 96513 48945 96559
rect 48991 96513 49069 96559
rect 49115 96513 49193 96559
rect 49239 96513 49317 96559
rect 49363 96513 49441 96559
rect 49487 96513 49565 96559
rect 49611 96513 49689 96559
rect 49735 96513 49813 96559
rect 49859 96513 49937 96559
rect 49983 96513 50061 96559
rect 50107 96513 50185 96559
rect 50231 96513 50309 96559
rect 50355 96513 50433 96559
rect 50479 96513 50557 96559
rect 50603 96513 50681 96559
rect 50727 96513 50805 96559
rect 50851 96513 50929 96559
rect 50975 96513 51053 96559
rect 51099 96513 51177 96559
rect 51223 96513 51301 96559
rect 51347 96513 51425 96559
rect 51471 96513 51549 96559
rect 51595 96513 51673 96559
rect 51719 96513 51797 96559
rect 51843 96513 51921 96559
rect 51967 96513 52045 96559
rect 52091 96513 52169 96559
rect 52215 96513 52293 96559
rect 52339 96513 52417 96559
rect 52463 96513 52541 96559
rect 52587 96513 52665 96559
rect 52711 96513 52789 96559
rect 52835 96513 52913 96559
rect 52959 96513 53037 96559
rect 53083 96513 53161 96559
rect 53207 96513 53285 96559
rect 53331 96513 53409 96559
rect 53455 96513 53533 96559
rect 53579 96513 53657 96559
rect 53703 96513 53781 96559
rect 53827 96513 53905 96559
rect 53951 96513 54029 96559
rect 54075 96513 54153 96559
rect 54199 96513 54277 96559
rect 54323 96513 54401 96559
rect 54447 96513 54525 96559
rect 54571 96513 54649 96559
rect 54695 96513 54773 96559
rect 54819 96513 54897 96559
rect 54943 96513 55021 96559
rect 55067 96513 55145 96559
rect 55191 96513 55269 96559
rect 55315 96513 55393 96559
rect 55439 96513 55517 96559
rect 55563 96513 55641 96559
rect 55687 96513 55765 96559
rect 55811 96513 55889 96559
rect 55935 96513 56013 96559
rect 56059 96513 56137 96559
rect 56183 96513 56261 96559
rect 56307 96513 56385 96559
rect 56431 96513 56509 96559
rect 56555 96513 56633 96559
rect 56679 96513 56757 96559
rect 56803 96513 56881 96559
rect 56927 96513 57005 96559
rect 57051 96513 57129 96559
rect 57175 96513 57253 96559
rect 57299 96513 57377 96559
rect 57423 96513 57501 96559
rect 57547 96513 57625 96559
rect 57671 96513 57749 96559
rect 57795 96513 57873 96559
rect 57919 96513 57997 96559
rect 58043 96513 58121 96559
rect 58167 96513 58245 96559
rect 58291 96513 58369 96559
rect 58415 96513 58493 96559
rect 58539 96513 58617 96559
rect 58663 96513 58741 96559
rect 58787 96513 58865 96559
rect 58911 96513 58989 96559
rect 59035 96513 59113 96559
rect 59159 96513 59237 96559
rect 59283 96513 59361 96559
rect 59407 96513 59485 96559
rect 59531 96513 59609 96559
rect 59655 96513 59733 96559
rect 59779 96513 59857 96559
rect 59903 96513 59981 96559
rect 60027 96513 60105 96559
rect 60151 96513 60229 96559
rect 60275 96513 60353 96559
rect 60399 96513 60477 96559
rect 60523 96513 60601 96559
rect 60647 96513 60725 96559
rect 60771 96513 60849 96559
rect 60895 96513 60973 96559
rect 61019 96513 61097 96559
rect 61143 96513 61221 96559
rect 61267 96513 61345 96559
rect 61391 96513 61469 96559
rect 61515 96513 61593 96559
rect 61639 96513 61717 96559
rect 61763 96513 61841 96559
rect 61887 96513 61965 96559
rect 62011 96513 62089 96559
rect 62135 96513 62213 96559
rect 62259 96513 62337 96559
rect 62383 96513 62461 96559
rect 62507 96513 62585 96559
rect 62631 96513 62709 96559
rect 62755 96513 62833 96559
rect 62879 96513 62957 96559
rect 63003 96513 63081 96559
rect 63127 96513 63205 96559
rect 63251 96513 63329 96559
rect 63375 96513 63453 96559
rect 63499 96513 63577 96559
rect 63623 96513 63701 96559
rect 63747 96513 63825 96559
rect 63871 96513 63949 96559
rect 63995 96513 64073 96559
rect 64119 96513 64197 96559
rect 64243 96513 64321 96559
rect 64367 96513 64445 96559
rect 64491 96513 64569 96559
rect 64615 96513 64693 96559
rect 64739 96513 64817 96559
rect 64863 96513 64941 96559
rect 64987 96513 65065 96559
rect 65111 96513 65189 96559
rect 65235 96513 65313 96559
rect 65359 96513 65437 96559
rect 65483 96513 65561 96559
rect 65607 96513 65685 96559
rect 65731 96513 65809 96559
rect 65855 96513 65933 96559
rect 65979 96513 66057 96559
rect 66103 96513 66181 96559
rect 66227 96513 66305 96559
rect 66351 96513 66429 96559
rect 66475 96513 66553 96559
rect 66599 96513 66677 96559
rect 66723 96513 66801 96559
rect 66847 96513 66925 96559
rect 66971 96513 67049 96559
rect 67095 96513 67173 96559
rect 67219 96513 67297 96559
rect 67343 96513 67421 96559
rect 67467 96513 67545 96559
rect 67591 96513 67669 96559
rect 67715 96513 67793 96559
rect 67839 96513 67917 96559
rect 67963 96513 68041 96559
rect 68087 96513 68165 96559
rect 68211 96513 68289 96559
rect 68335 96513 68413 96559
rect 68459 96513 68537 96559
rect 68583 96513 68661 96559
rect 68707 96513 68785 96559
rect 68831 96513 68909 96559
rect 68955 96513 69033 96559
rect 69079 96513 69157 96559
rect 69203 96513 69281 96559
rect 69327 96513 69405 96559
rect 69451 96513 69529 96559
rect 69575 96513 69653 96559
rect 69699 96513 69777 96559
rect 69823 96513 69901 96559
rect 69947 96513 70025 96559
rect 70071 96513 70149 96559
rect 70195 96513 70273 96559
rect 70319 96513 70397 96559
rect 70443 96513 70521 96559
rect 70567 96513 70645 96559
rect 70691 96513 70769 96559
rect 70815 96513 70893 96559
rect 70939 96513 71017 96559
rect 71063 96513 71141 96559
rect 71187 96513 71265 96559
rect 71311 96513 71389 96559
rect 71435 96513 71513 96559
rect 71559 96513 71637 96559
rect 71683 96513 71761 96559
rect 71807 96513 71885 96559
rect 71931 96513 72009 96559
rect 72055 96513 72133 96559
rect 72179 96513 72257 96559
rect 72303 96513 72381 96559
rect 72427 96513 72505 96559
rect 72551 96513 72629 96559
rect 72675 96513 72753 96559
rect 72799 96513 72877 96559
rect 72923 96513 73001 96559
rect 73047 96513 73125 96559
rect 73171 96513 73249 96559
rect 73295 96513 73373 96559
rect 73419 96513 73497 96559
rect 73543 96513 73621 96559
rect 73667 96513 73745 96559
rect 73791 96513 73869 96559
rect 73915 96513 73993 96559
rect 74039 96513 74117 96559
rect 74163 96513 74241 96559
rect 74287 96513 74365 96559
rect 74411 96513 74489 96559
rect 74535 96513 74613 96559
rect 74659 96513 74737 96559
rect 74783 96513 74861 96559
rect 74907 96513 74985 96559
rect 75031 96513 75109 96559
rect 75155 96513 75233 96559
rect 75279 96513 75357 96559
rect 75403 96513 75481 96559
rect 75527 96513 75605 96559
rect 75651 96513 75729 96559
rect 75775 96513 75853 96559
rect 75899 96513 75977 96559
rect 76023 96513 76101 96559
rect 76147 96513 76225 96559
rect 76271 96513 76349 96559
rect 76395 96513 76473 96559
rect 76519 96513 76597 96559
rect 76643 96513 76721 96559
rect 76767 96513 76845 96559
rect 76891 96513 76969 96559
rect 77015 96513 77093 96559
rect 77139 96513 77217 96559
rect 77263 96513 77341 96559
rect 77387 96513 77465 96559
rect 77511 96513 77589 96559
rect 77635 96513 77713 96559
rect 77759 96513 77837 96559
rect 77883 96513 77961 96559
rect 78007 96513 78085 96559
rect 78131 96513 78209 96559
rect 78255 96513 78333 96559
rect 78379 96513 78457 96559
rect 78503 96513 78581 96559
rect 78627 96513 78705 96559
rect 78751 96513 78829 96559
rect 78875 96513 78953 96559
rect 78999 96513 79077 96559
rect 79123 96513 79201 96559
rect 79247 96513 79325 96559
rect 79371 96513 79449 96559
rect 79495 96513 79573 96559
rect 79619 96513 79697 96559
rect 79743 96513 79821 96559
rect 79867 96513 79945 96559
rect 79991 96513 80069 96559
rect 80115 96513 80193 96559
rect 80239 96513 80317 96559
rect 80363 96513 80441 96559
rect 80487 96513 80565 96559
rect 80611 96513 80689 96559
rect 80735 96513 80813 96559
rect 80859 96513 80937 96559
rect 80983 96513 81061 96559
rect 81107 96513 81185 96559
rect 81231 96513 81309 96559
rect 81355 96513 81433 96559
rect 81479 96513 81557 96559
rect 81603 96513 81681 96559
rect 81727 96513 81805 96559
rect 81851 96513 81929 96559
rect 81975 96513 82053 96559
rect 82099 96513 82177 96559
rect 82223 96513 82301 96559
rect 82347 96513 82425 96559
rect 82471 96513 82549 96559
rect 82595 96513 82673 96559
rect 82719 96513 82797 96559
rect 82843 96513 82921 96559
rect 82967 96513 83045 96559
rect 83091 96513 83169 96559
rect 83215 96513 83293 96559
rect 83339 96513 83417 96559
rect 83463 96513 83541 96559
rect 83587 96513 83665 96559
rect 83711 96513 83789 96559
rect 83835 96513 83913 96559
rect 83959 96513 84037 96559
rect 84083 96513 84161 96559
rect 84207 96513 84285 96559
rect 84331 96513 84409 96559
rect 84455 96513 84533 96559
rect 84579 96513 84657 96559
rect 84703 96513 84781 96559
rect 84827 96513 84905 96559
rect 84951 96513 85029 96559
rect 85075 96513 85153 96559
rect 85199 96513 85277 96559
rect 85323 96513 85401 96559
rect 85447 96513 85525 96559
rect 85571 96513 85649 96559
rect 85695 96513 85706 96559
rect 0 96435 85706 96513
rect 0 96389 89 96435
rect 135 96389 213 96435
rect 259 96389 337 96435
rect 383 96389 461 96435
rect 507 96389 585 96435
rect 631 96389 709 96435
rect 755 96389 833 96435
rect 879 96389 957 96435
rect 1003 96389 1081 96435
rect 1127 96389 1205 96435
rect 1251 96389 1329 96435
rect 1375 96389 1453 96435
rect 1499 96389 1577 96435
rect 1623 96389 1701 96435
rect 1747 96389 1825 96435
rect 1871 96389 1949 96435
rect 1995 96389 2073 96435
rect 2119 96389 2197 96435
rect 2243 96389 2321 96435
rect 2367 96389 2445 96435
rect 2491 96389 2569 96435
rect 2615 96389 2693 96435
rect 2739 96389 2817 96435
rect 2863 96389 2941 96435
rect 2987 96389 3065 96435
rect 3111 96389 3189 96435
rect 3235 96389 3313 96435
rect 3359 96389 3437 96435
rect 3483 96389 3561 96435
rect 3607 96389 3685 96435
rect 3731 96389 3809 96435
rect 3855 96389 3933 96435
rect 3979 96389 4057 96435
rect 4103 96389 4181 96435
rect 4227 96389 4305 96435
rect 4351 96389 4429 96435
rect 4475 96389 4553 96435
rect 4599 96389 4677 96435
rect 4723 96389 4801 96435
rect 4847 96389 4925 96435
rect 4971 96389 5049 96435
rect 5095 96389 5173 96435
rect 5219 96389 5297 96435
rect 5343 96389 5421 96435
rect 5467 96389 5545 96435
rect 5591 96389 5669 96435
rect 5715 96389 5793 96435
rect 5839 96389 5917 96435
rect 5963 96389 6041 96435
rect 6087 96389 6165 96435
rect 6211 96389 6289 96435
rect 6335 96389 6413 96435
rect 6459 96389 6537 96435
rect 6583 96389 6661 96435
rect 6707 96389 6785 96435
rect 6831 96389 6909 96435
rect 6955 96389 7033 96435
rect 7079 96389 7157 96435
rect 7203 96389 7281 96435
rect 7327 96389 7405 96435
rect 7451 96389 7529 96435
rect 7575 96389 7653 96435
rect 7699 96389 7777 96435
rect 7823 96389 7901 96435
rect 7947 96389 8025 96435
rect 8071 96389 8149 96435
rect 8195 96389 8273 96435
rect 8319 96389 8397 96435
rect 8443 96389 8521 96435
rect 8567 96389 8645 96435
rect 8691 96389 8769 96435
rect 8815 96389 8893 96435
rect 8939 96389 9017 96435
rect 9063 96389 9141 96435
rect 9187 96389 9265 96435
rect 9311 96389 9389 96435
rect 9435 96389 9513 96435
rect 9559 96389 9637 96435
rect 9683 96389 9761 96435
rect 9807 96389 9885 96435
rect 9931 96389 10009 96435
rect 10055 96389 10133 96435
rect 10179 96389 10257 96435
rect 10303 96389 10381 96435
rect 10427 96389 10505 96435
rect 10551 96389 10629 96435
rect 10675 96389 10753 96435
rect 10799 96389 10877 96435
rect 10923 96389 11001 96435
rect 11047 96389 11125 96435
rect 11171 96389 11249 96435
rect 11295 96389 11373 96435
rect 11419 96389 11497 96435
rect 11543 96389 11621 96435
rect 11667 96389 11745 96435
rect 11791 96389 11869 96435
rect 11915 96389 11993 96435
rect 12039 96389 12117 96435
rect 12163 96389 12241 96435
rect 12287 96389 12365 96435
rect 12411 96389 12489 96435
rect 12535 96389 12613 96435
rect 12659 96389 12737 96435
rect 12783 96389 12861 96435
rect 12907 96389 12985 96435
rect 13031 96389 13109 96435
rect 13155 96389 13233 96435
rect 13279 96389 13357 96435
rect 13403 96389 13481 96435
rect 13527 96389 13605 96435
rect 13651 96389 13729 96435
rect 13775 96389 13853 96435
rect 13899 96389 13977 96435
rect 14023 96389 14101 96435
rect 14147 96389 14225 96435
rect 14271 96389 14349 96435
rect 14395 96389 14473 96435
rect 14519 96389 14597 96435
rect 14643 96389 14721 96435
rect 14767 96389 14845 96435
rect 14891 96389 14969 96435
rect 15015 96389 15093 96435
rect 15139 96389 15217 96435
rect 15263 96389 15341 96435
rect 15387 96389 15465 96435
rect 15511 96389 15589 96435
rect 15635 96389 15713 96435
rect 15759 96389 15837 96435
rect 15883 96389 15961 96435
rect 16007 96389 16085 96435
rect 16131 96389 16209 96435
rect 16255 96389 16333 96435
rect 16379 96389 16457 96435
rect 16503 96389 16581 96435
rect 16627 96389 16705 96435
rect 16751 96389 16829 96435
rect 16875 96389 16953 96435
rect 16999 96389 17077 96435
rect 17123 96389 17201 96435
rect 17247 96389 17325 96435
rect 17371 96389 17449 96435
rect 17495 96389 17573 96435
rect 17619 96389 17697 96435
rect 17743 96389 17821 96435
rect 17867 96389 17945 96435
rect 17991 96389 18069 96435
rect 18115 96389 18193 96435
rect 18239 96389 18317 96435
rect 18363 96389 18441 96435
rect 18487 96389 18565 96435
rect 18611 96389 18689 96435
rect 18735 96389 18813 96435
rect 18859 96389 18937 96435
rect 18983 96389 19061 96435
rect 19107 96389 19185 96435
rect 19231 96389 19309 96435
rect 19355 96389 19433 96435
rect 19479 96389 19557 96435
rect 19603 96389 19681 96435
rect 19727 96389 19805 96435
rect 19851 96389 19929 96435
rect 19975 96389 20053 96435
rect 20099 96389 20177 96435
rect 20223 96389 20301 96435
rect 20347 96389 20425 96435
rect 20471 96389 20549 96435
rect 20595 96389 20673 96435
rect 20719 96389 20797 96435
rect 20843 96389 20921 96435
rect 20967 96389 21045 96435
rect 21091 96389 21169 96435
rect 21215 96389 21293 96435
rect 21339 96389 21417 96435
rect 21463 96389 21541 96435
rect 21587 96389 21665 96435
rect 21711 96389 21789 96435
rect 21835 96389 21913 96435
rect 21959 96389 22037 96435
rect 22083 96389 22161 96435
rect 22207 96389 22285 96435
rect 22331 96389 22409 96435
rect 22455 96389 22533 96435
rect 22579 96389 22657 96435
rect 22703 96389 22781 96435
rect 22827 96389 22905 96435
rect 22951 96389 23029 96435
rect 23075 96389 23153 96435
rect 23199 96389 23277 96435
rect 23323 96389 23401 96435
rect 23447 96389 23525 96435
rect 23571 96389 23649 96435
rect 23695 96389 23773 96435
rect 23819 96389 23897 96435
rect 23943 96389 24021 96435
rect 24067 96389 24145 96435
rect 24191 96389 24269 96435
rect 24315 96389 24393 96435
rect 24439 96389 24517 96435
rect 24563 96389 24641 96435
rect 24687 96389 24765 96435
rect 24811 96389 24889 96435
rect 24935 96389 25013 96435
rect 25059 96389 25137 96435
rect 25183 96389 25261 96435
rect 25307 96389 25385 96435
rect 25431 96389 25509 96435
rect 25555 96389 25633 96435
rect 25679 96389 25757 96435
rect 25803 96389 25881 96435
rect 25927 96389 26005 96435
rect 26051 96389 26129 96435
rect 26175 96389 26253 96435
rect 26299 96389 26377 96435
rect 26423 96389 26501 96435
rect 26547 96389 26625 96435
rect 26671 96389 26749 96435
rect 26795 96389 26873 96435
rect 26919 96389 26997 96435
rect 27043 96389 27121 96435
rect 27167 96389 27245 96435
rect 27291 96389 27369 96435
rect 27415 96389 27493 96435
rect 27539 96389 27617 96435
rect 27663 96389 27741 96435
rect 27787 96389 27865 96435
rect 27911 96389 27989 96435
rect 28035 96389 28113 96435
rect 28159 96389 28237 96435
rect 28283 96389 28361 96435
rect 28407 96389 28485 96435
rect 28531 96389 28609 96435
rect 28655 96389 28733 96435
rect 28779 96389 28857 96435
rect 28903 96389 28981 96435
rect 29027 96389 29105 96435
rect 29151 96389 29229 96435
rect 29275 96389 29353 96435
rect 29399 96389 29477 96435
rect 29523 96389 29601 96435
rect 29647 96389 29725 96435
rect 29771 96389 29849 96435
rect 29895 96389 29973 96435
rect 30019 96389 30097 96435
rect 30143 96389 30221 96435
rect 30267 96389 30345 96435
rect 30391 96389 30469 96435
rect 30515 96389 30593 96435
rect 30639 96389 30717 96435
rect 30763 96389 30841 96435
rect 30887 96389 30965 96435
rect 31011 96389 31089 96435
rect 31135 96389 31213 96435
rect 31259 96389 31337 96435
rect 31383 96389 31461 96435
rect 31507 96389 31585 96435
rect 31631 96389 31709 96435
rect 31755 96389 31833 96435
rect 31879 96389 31957 96435
rect 32003 96389 32081 96435
rect 32127 96389 32205 96435
rect 32251 96389 32329 96435
rect 32375 96389 32453 96435
rect 32499 96389 32577 96435
rect 32623 96389 32701 96435
rect 32747 96389 32825 96435
rect 32871 96389 32949 96435
rect 32995 96389 33073 96435
rect 33119 96389 33197 96435
rect 33243 96389 33321 96435
rect 33367 96389 33445 96435
rect 33491 96389 33569 96435
rect 33615 96389 33693 96435
rect 33739 96389 33817 96435
rect 33863 96389 33941 96435
rect 33987 96389 34065 96435
rect 34111 96389 34189 96435
rect 34235 96389 34313 96435
rect 34359 96389 34437 96435
rect 34483 96389 34561 96435
rect 34607 96389 34685 96435
rect 34731 96389 34809 96435
rect 34855 96389 34933 96435
rect 34979 96389 35057 96435
rect 35103 96389 35181 96435
rect 35227 96389 35305 96435
rect 35351 96389 35429 96435
rect 35475 96389 35553 96435
rect 35599 96389 35677 96435
rect 35723 96389 35801 96435
rect 35847 96389 35925 96435
rect 35971 96389 36049 96435
rect 36095 96389 36173 96435
rect 36219 96389 36297 96435
rect 36343 96389 36421 96435
rect 36467 96389 36545 96435
rect 36591 96389 36669 96435
rect 36715 96389 36793 96435
rect 36839 96389 36917 96435
rect 36963 96389 37041 96435
rect 37087 96389 37165 96435
rect 37211 96389 37289 96435
rect 37335 96389 37413 96435
rect 37459 96389 37537 96435
rect 37583 96389 37661 96435
rect 37707 96389 37785 96435
rect 37831 96389 37909 96435
rect 37955 96389 38033 96435
rect 38079 96389 38157 96435
rect 38203 96389 38281 96435
rect 38327 96389 38405 96435
rect 38451 96389 38529 96435
rect 38575 96389 38653 96435
rect 38699 96389 38777 96435
rect 38823 96389 38901 96435
rect 38947 96389 39025 96435
rect 39071 96389 39149 96435
rect 39195 96389 39273 96435
rect 39319 96389 39397 96435
rect 39443 96389 39521 96435
rect 39567 96389 39645 96435
rect 39691 96389 39769 96435
rect 39815 96389 39893 96435
rect 39939 96389 40017 96435
rect 40063 96389 40141 96435
rect 40187 96389 40265 96435
rect 40311 96389 40389 96435
rect 40435 96389 40513 96435
rect 40559 96389 40637 96435
rect 40683 96389 40761 96435
rect 40807 96389 40885 96435
rect 40931 96389 41009 96435
rect 41055 96389 41133 96435
rect 41179 96389 41257 96435
rect 41303 96389 41381 96435
rect 41427 96389 41505 96435
rect 41551 96389 41629 96435
rect 41675 96389 41753 96435
rect 41799 96389 41877 96435
rect 41923 96389 42001 96435
rect 42047 96389 42125 96435
rect 42171 96389 42249 96435
rect 42295 96389 42373 96435
rect 42419 96389 42497 96435
rect 42543 96389 42621 96435
rect 42667 96389 42745 96435
rect 42791 96389 42869 96435
rect 42915 96389 42993 96435
rect 43039 96389 43117 96435
rect 43163 96389 43241 96435
rect 43287 96389 43365 96435
rect 43411 96389 43489 96435
rect 43535 96389 43613 96435
rect 43659 96389 43737 96435
rect 43783 96389 43861 96435
rect 43907 96389 43985 96435
rect 44031 96389 44109 96435
rect 44155 96389 44233 96435
rect 44279 96389 44357 96435
rect 44403 96389 44481 96435
rect 44527 96389 44605 96435
rect 44651 96389 44729 96435
rect 44775 96389 44853 96435
rect 44899 96389 44977 96435
rect 45023 96389 45101 96435
rect 45147 96389 45225 96435
rect 45271 96389 45349 96435
rect 45395 96389 45473 96435
rect 45519 96389 45597 96435
rect 45643 96389 45721 96435
rect 45767 96389 45845 96435
rect 45891 96389 45969 96435
rect 46015 96389 46093 96435
rect 46139 96389 46217 96435
rect 46263 96389 46341 96435
rect 46387 96389 46465 96435
rect 46511 96389 46589 96435
rect 46635 96389 46713 96435
rect 46759 96389 46837 96435
rect 46883 96389 46961 96435
rect 47007 96389 47085 96435
rect 47131 96389 47209 96435
rect 47255 96389 47333 96435
rect 47379 96389 47457 96435
rect 47503 96389 47581 96435
rect 47627 96389 47705 96435
rect 47751 96389 47829 96435
rect 47875 96389 47953 96435
rect 47999 96389 48077 96435
rect 48123 96389 48201 96435
rect 48247 96389 48325 96435
rect 48371 96389 48449 96435
rect 48495 96389 48573 96435
rect 48619 96389 48697 96435
rect 48743 96389 48821 96435
rect 48867 96389 48945 96435
rect 48991 96389 49069 96435
rect 49115 96389 49193 96435
rect 49239 96389 49317 96435
rect 49363 96389 49441 96435
rect 49487 96389 49565 96435
rect 49611 96389 49689 96435
rect 49735 96389 49813 96435
rect 49859 96389 49937 96435
rect 49983 96389 50061 96435
rect 50107 96389 50185 96435
rect 50231 96389 50309 96435
rect 50355 96389 50433 96435
rect 50479 96389 50557 96435
rect 50603 96389 50681 96435
rect 50727 96389 50805 96435
rect 50851 96389 50929 96435
rect 50975 96389 51053 96435
rect 51099 96389 51177 96435
rect 51223 96389 51301 96435
rect 51347 96389 51425 96435
rect 51471 96389 51549 96435
rect 51595 96389 51673 96435
rect 51719 96389 51797 96435
rect 51843 96389 51921 96435
rect 51967 96389 52045 96435
rect 52091 96389 52169 96435
rect 52215 96389 52293 96435
rect 52339 96389 52417 96435
rect 52463 96389 52541 96435
rect 52587 96389 52665 96435
rect 52711 96389 52789 96435
rect 52835 96389 52913 96435
rect 52959 96389 53037 96435
rect 53083 96389 53161 96435
rect 53207 96389 53285 96435
rect 53331 96389 53409 96435
rect 53455 96389 53533 96435
rect 53579 96389 53657 96435
rect 53703 96389 53781 96435
rect 53827 96389 53905 96435
rect 53951 96389 54029 96435
rect 54075 96389 54153 96435
rect 54199 96389 54277 96435
rect 54323 96389 54401 96435
rect 54447 96389 54525 96435
rect 54571 96389 54649 96435
rect 54695 96389 54773 96435
rect 54819 96389 54897 96435
rect 54943 96389 55021 96435
rect 55067 96389 55145 96435
rect 55191 96389 55269 96435
rect 55315 96389 55393 96435
rect 55439 96389 55517 96435
rect 55563 96389 55641 96435
rect 55687 96389 55765 96435
rect 55811 96389 55889 96435
rect 55935 96389 56013 96435
rect 56059 96389 56137 96435
rect 56183 96389 56261 96435
rect 56307 96389 56385 96435
rect 56431 96389 56509 96435
rect 56555 96389 56633 96435
rect 56679 96389 56757 96435
rect 56803 96389 56881 96435
rect 56927 96389 57005 96435
rect 57051 96389 57129 96435
rect 57175 96389 57253 96435
rect 57299 96389 57377 96435
rect 57423 96389 57501 96435
rect 57547 96389 57625 96435
rect 57671 96389 57749 96435
rect 57795 96389 57873 96435
rect 57919 96389 57997 96435
rect 58043 96389 58121 96435
rect 58167 96389 58245 96435
rect 58291 96389 58369 96435
rect 58415 96389 58493 96435
rect 58539 96389 58617 96435
rect 58663 96389 58741 96435
rect 58787 96389 58865 96435
rect 58911 96389 58989 96435
rect 59035 96389 59113 96435
rect 59159 96389 59237 96435
rect 59283 96389 59361 96435
rect 59407 96389 59485 96435
rect 59531 96389 59609 96435
rect 59655 96389 59733 96435
rect 59779 96389 59857 96435
rect 59903 96389 59981 96435
rect 60027 96389 60105 96435
rect 60151 96389 60229 96435
rect 60275 96389 60353 96435
rect 60399 96389 60477 96435
rect 60523 96389 60601 96435
rect 60647 96389 60725 96435
rect 60771 96389 60849 96435
rect 60895 96389 60973 96435
rect 61019 96389 61097 96435
rect 61143 96389 61221 96435
rect 61267 96389 61345 96435
rect 61391 96389 61469 96435
rect 61515 96389 61593 96435
rect 61639 96389 61717 96435
rect 61763 96389 61841 96435
rect 61887 96389 61965 96435
rect 62011 96389 62089 96435
rect 62135 96389 62213 96435
rect 62259 96389 62337 96435
rect 62383 96389 62461 96435
rect 62507 96389 62585 96435
rect 62631 96389 62709 96435
rect 62755 96389 62833 96435
rect 62879 96389 62957 96435
rect 63003 96389 63081 96435
rect 63127 96389 63205 96435
rect 63251 96389 63329 96435
rect 63375 96389 63453 96435
rect 63499 96389 63577 96435
rect 63623 96389 63701 96435
rect 63747 96389 63825 96435
rect 63871 96389 63949 96435
rect 63995 96389 64073 96435
rect 64119 96389 64197 96435
rect 64243 96389 64321 96435
rect 64367 96389 64445 96435
rect 64491 96389 64569 96435
rect 64615 96389 64693 96435
rect 64739 96389 64817 96435
rect 64863 96389 64941 96435
rect 64987 96389 65065 96435
rect 65111 96389 65189 96435
rect 65235 96389 65313 96435
rect 65359 96389 65437 96435
rect 65483 96389 65561 96435
rect 65607 96389 65685 96435
rect 65731 96389 65809 96435
rect 65855 96389 65933 96435
rect 65979 96389 66057 96435
rect 66103 96389 66181 96435
rect 66227 96389 66305 96435
rect 66351 96389 66429 96435
rect 66475 96389 66553 96435
rect 66599 96389 66677 96435
rect 66723 96389 66801 96435
rect 66847 96389 66925 96435
rect 66971 96389 67049 96435
rect 67095 96389 67173 96435
rect 67219 96389 67297 96435
rect 67343 96389 67421 96435
rect 67467 96389 67545 96435
rect 67591 96389 67669 96435
rect 67715 96389 67793 96435
rect 67839 96389 67917 96435
rect 67963 96389 68041 96435
rect 68087 96389 68165 96435
rect 68211 96389 68289 96435
rect 68335 96389 68413 96435
rect 68459 96389 68537 96435
rect 68583 96389 68661 96435
rect 68707 96389 68785 96435
rect 68831 96389 68909 96435
rect 68955 96389 69033 96435
rect 69079 96389 69157 96435
rect 69203 96389 69281 96435
rect 69327 96389 69405 96435
rect 69451 96389 69529 96435
rect 69575 96389 69653 96435
rect 69699 96389 69777 96435
rect 69823 96389 69901 96435
rect 69947 96389 70025 96435
rect 70071 96389 70149 96435
rect 70195 96389 70273 96435
rect 70319 96389 70397 96435
rect 70443 96389 70521 96435
rect 70567 96389 70645 96435
rect 70691 96389 70769 96435
rect 70815 96389 70893 96435
rect 70939 96389 71017 96435
rect 71063 96389 71141 96435
rect 71187 96389 71265 96435
rect 71311 96389 71389 96435
rect 71435 96389 71513 96435
rect 71559 96389 71637 96435
rect 71683 96389 71761 96435
rect 71807 96389 71885 96435
rect 71931 96389 72009 96435
rect 72055 96389 72133 96435
rect 72179 96389 72257 96435
rect 72303 96389 72381 96435
rect 72427 96389 72505 96435
rect 72551 96389 72629 96435
rect 72675 96389 72753 96435
rect 72799 96389 72877 96435
rect 72923 96389 73001 96435
rect 73047 96389 73125 96435
rect 73171 96389 73249 96435
rect 73295 96389 73373 96435
rect 73419 96389 73497 96435
rect 73543 96389 73621 96435
rect 73667 96389 73745 96435
rect 73791 96389 73869 96435
rect 73915 96389 73993 96435
rect 74039 96389 74117 96435
rect 74163 96389 74241 96435
rect 74287 96389 74365 96435
rect 74411 96389 74489 96435
rect 74535 96389 74613 96435
rect 74659 96389 74737 96435
rect 74783 96389 74861 96435
rect 74907 96389 74985 96435
rect 75031 96389 75109 96435
rect 75155 96389 75233 96435
rect 75279 96389 75357 96435
rect 75403 96389 75481 96435
rect 75527 96389 75605 96435
rect 75651 96389 75729 96435
rect 75775 96389 75853 96435
rect 75899 96389 75977 96435
rect 76023 96389 76101 96435
rect 76147 96389 76225 96435
rect 76271 96389 76349 96435
rect 76395 96389 76473 96435
rect 76519 96389 76597 96435
rect 76643 96389 76721 96435
rect 76767 96389 76845 96435
rect 76891 96389 76969 96435
rect 77015 96389 77093 96435
rect 77139 96389 77217 96435
rect 77263 96389 77341 96435
rect 77387 96389 77465 96435
rect 77511 96389 77589 96435
rect 77635 96389 77713 96435
rect 77759 96389 77837 96435
rect 77883 96389 77961 96435
rect 78007 96389 78085 96435
rect 78131 96389 78209 96435
rect 78255 96389 78333 96435
rect 78379 96389 78457 96435
rect 78503 96389 78581 96435
rect 78627 96389 78705 96435
rect 78751 96389 78829 96435
rect 78875 96389 78953 96435
rect 78999 96389 79077 96435
rect 79123 96389 79201 96435
rect 79247 96389 79325 96435
rect 79371 96389 79449 96435
rect 79495 96389 79573 96435
rect 79619 96389 79697 96435
rect 79743 96389 79821 96435
rect 79867 96389 79945 96435
rect 79991 96389 80069 96435
rect 80115 96389 80193 96435
rect 80239 96389 80317 96435
rect 80363 96389 80441 96435
rect 80487 96389 80565 96435
rect 80611 96389 80689 96435
rect 80735 96389 80813 96435
rect 80859 96389 80937 96435
rect 80983 96389 81061 96435
rect 81107 96389 81185 96435
rect 81231 96389 81309 96435
rect 81355 96389 81433 96435
rect 81479 96389 81557 96435
rect 81603 96389 81681 96435
rect 81727 96389 81805 96435
rect 81851 96389 81929 96435
rect 81975 96389 82053 96435
rect 82099 96389 82177 96435
rect 82223 96389 82301 96435
rect 82347 96389 82425 96435
rect 82471 96389 82549 96435
rect 82595 96389 82673 96435
rect 82719 96389 82797 96435
rect 82843 96389 82921 96435
rect 82967 96389 83045 96435
rect 83091 96389 83169 96435
rect 83215 96389 83293 96435
rect 83339 96389 83417 96435
rect 83463 96389 83541 96435
rect 83587 96389 83665 96435
rect 83711 96389 83789 96435
rect 83835 96389 83913 96435
rect 83959 96389 84037 96435
rect 84083 96389 84161 96435
rect 84207 96389 84285 96435
rect 84331 96389 84409 96435
rect 84455 96389 84533 96435
rect 84579 96389 84657 96435
rect 84703 96389 84781 96435
rect 84827 96389 84905 96435
rect 84951 96389 85029 96435
rect 85075 96389 85153 96435
rect 85199 96389 85277 96435
rect 85323 96389 85401 96435
rect 85447 96389 85525 96435
rect 85571 96389 85649 96435
rect 85695 96389 85706 96435
rect 0 96311 85706 96389
rect 0 96265 89 96311
rect 135 96265 213 96311
rect 259 96265 337 96311
rect 383 96265 461 96311
rect 507 96265 585 96311
rect 631 96265 709 96311
rect 755 96265 833 96311
rect 879 96265 957 96311
rect 1003 96265 1081 96311
rect 1127 96265 1205 96311
rect 1251 96265 1329 96311
rect 1375 96265 1453 96311
rect 1499 96265 1577 96311
rect 1623 96265 1701 96311
rect 1747 96265 1825 96311
rect 1871 96265 1949 96311
rect 1995 96265 2073 96311
rect 2119 96265 2197 96311
rect 2243 96265 2321 96311
rect 2367 96265 2445 96311
rect 2491 96265 2569 96311
rect 2615 96265 2693 96311
rect 2739 96265 2817 96311
rect 2863 96265 2941 96311
rect 2987 96265 3065 96311
rect 3111 96265 3189 96311
rect 3235 96265 3313 96311
rect 3359 96265 3437 96311
rect 3483 96265 3561 96311
rect 3607 96265 3685 96311
rect 3731 96265 3809 96311
rect 3855 96265 3933 96311
rect 3979 96265 4057 96311
rect 4103 96265 4181 96311
rect 4227 96265 4305 96311
rect 4351 96265 4429 96311
rect 4475 96265 4553 96311
rect 4599 96265 4677 96311
rect 4723 96265 4801 96311
rect 4847 96265 4925 96311
rect 4971 96265 5049 96311
rect 5095 96265 5173 96311
rect 5219 96265 5297 96311
rect 5343 96265 5421 96311
rect 5467 96265 5545 96311
rect 5591 96265 5669 96311
rect 5715 96265 5793 96311
rect 5839 96265 5917 96311
rect 5963 96265 6041 96311
rect 6087 96265 6165 96311
rect 6211 96265 6289 96311
rect 6335 96265 6413 96311
rect 6459 96265 6537 96311
rect 6583 96265 6661 96311
rect 6707 96265 6785 96311
rect 6831 96265 6909 96311
rect 6955 96265 7033 96311
rect 7079 96265 7157 96311
rect 7203 96265 7281 96311
rect 7327 96265 7405 96311
rect 7451 96265 7529 96311
rect 7575 96265 7653 96311
rect 7699 96265 7777 96311
rect 7823 96265 7901 96311
rect 7947 96265 8025 96311
rect 8071 96265 8149 96311
rect 8195 96265 8273 96311
rect 8319 96265 8397 96311
rect 8443 96265 8521 96311
rect 8567 96265 8645 96311
rect 8691 96265 8769 96311
rect 8815 96265 8893 96311
rect 8939 96265 9017 96311
rect 9063 96265 9141 96311
rect 9187 96265 9265 96311
rect 9311 96265 9389 96311
rect 9435 96265 9513 96311
rect 9559 96265 9637 96311
rect 9683 96265 9761 96311
rect 9807 96265 9885 96311
rect 9931 96265 10009 96311
rect 10055 96265 10133 96311
rect 10179 96265 10257 96311
rect 10303 96265 10381 96311
rect 10427 96265 10505 96311
rect 10551 96265 10629 96311
rect 10675 96265 10753 96311
rect 10799 96265 10877 96311
rect 10923 96265 11001 96311
rect 11047 96265 11125 96311
rect 11171 96265 11249 96311
rect 11295 96265 11373 96311
rect 11419 96265 11497 96311
rect 11543 96265 11621 96311
rect 11667 96265 11745 96311
rect 11791 96265 11869 96311
rect 11915 96265 11993 96311
rect 12039 96265 12117 96311
rect 12163 96265 12241 96311
rect 12287 96265 12365 96311
rect 12411 96265 12489 96311
rect 12535 96265 12613 96311
rect 12659 96265 12737 96311
rect 12783 96265 12861 96311
rect 12907 96265 12985 96311
rect 13031 96265 13109 96311
rect 13155 96265 13233 96311
rect 13279 96265 13357 96311
rect 13403 96265 13481 96311
rect 13527 96265 13605 96311
rect 13651 96265 13729 96311
rect 13775 96265 13853 96311
rect 13899 96265 13977 96311
rect 14023 96265 14101 96311
rect 14147 96265 14225 96311
rect 14271 96265 14349 96311
rect 14395 96265 14473 96311
rect 14519 96265 14597 96311
rect 14643 96265 14721 96311
rect 14767 96265 14845 96311
rect 14891 96265 14969 96311
rect 15015 96265 15093 96311
rect 15139 96265 15217 96311
rect 15263 96265 15341 96311
rect 15387 96265 15465 96311
rect 15511 96265 15589 96311
rect 15635 96265 15713 96311
rect 15759 96265 15837 96311
rect 15883 96265 15961 96311
rect 16007 96265 16085 96311
rect 16131 96265 16209 96311
rect 16255 96265 16333 96311
rect 16379 96265 16457 96311
rect 16503 96265 16581 96311
rect 16627 96265 16705 96311
rect 16751 96265 16829 96311
rect 16875 96265 16953 96311
rect 16999 96265 17077 96311
rect 17123 96265 17201 96311
rect 17247 96265 17325 96311
rect 17371 96265 17449 96311
rect 17495 96265 17573 96311
rect 17619 96265 17697 96311
rect 17743 96265 17821 96311
rect 17867 96265 17945 96311
rect 17991 96265 18069 96311
rect 18115 96265 18193 96311
rect 18239 96265 18317 96311
rect 18363 96265 18441 96311
rect 18487 96265 18565 96311
rect 18611 96265 18689 96311
rect 18735 96265 18813 96311
rect 18859 96265 18937 96311
rect 18983 96265 19061 96311
rect 19107 96265 19185 96311
rect 19231 96265 19309 96311
rect 19355 96265 19433 96311
rect 19479 96265 19557 96311
rect 19603 96265 19681 96311
rect 19727 96265 19805 96311
rect 19851 96265 19929 96311
rect 19975 96265 20053 96311
rect 20099 96265 20177 96311
rect 20223 96265 20301 96311
rect 20347 96265 20425 96311
rect 20471 96265 20549 96311
rect 20595 96265 20673 96311
rect 20719 96265 20797 96311
rect 20843 96265 20921 96311
rect 20967 96265 21045 96311
rect 21091 96265 21169 96311
rect 21215 96265 21293 96311
rect 21339 96265 21417 96311
rect 21463 96265 21541 96311
rect 21587 96265 21665 96311
rect 21711 96265 21789 96311
rect 21835 96265 21913 96311
rect 21959 96265 22037 96311
rect 22083 96265 22161 96311
rect 22207 96265 22285 96311
rect 22331 96265 22409 96311
rect 22455 96265 22533 96311
rect 22579 96265 22657 96311
rect 22703 96265 22781 96311
rect 22827 96265 22905 96311
rect 22951 96265 23029 96311
rect 23075 96265 23153 96311
rect 23199 96265 23277 96311
rect 23323 96265 23401 96311
rect 23447 96265 23525 96311
rect 23571 96265 23649 96311
rect 23695 96265 23773 96311
rect 23819 96265 23897 96311
rect 23943 96265 24021 96311
rect 24067 96265 24145 96311
rect 24191 96265 24269 96311
rect 24315 96265 24393 96311
rect 24439 96265 24517 96311
rect 24563 96265 24641 96311
rect 24687 96265 24765 96311
rect 24811 96265 24889 96311
rect 24935 96265 25013 96311
rect 25059 96265 25137 96311
rect 25183 96265 25261 96311
rect 25307 96265 25385 96311
rect 25431 96265 25509 96311
rect 25555 96265 25633 96311
rect 25679 96265 25757 96311
rect 25803 96265 25881 96311
rect 25927 96265 26005 96311
rect 26051 96265 26129 96311
rect 26175 96265 26253 96311
rect 26299 96265 26377 96311
rect 26423 96265 26501 96311
rect 26547 96265 26625 96311
rect 26671 96265 26749 96311
rect 26795 96265 26873 96311
rect 26919 96265 26997 96311
rect 27043 96265 27121 96311
rect 27167 96265 27245 96311
rect 27291 96265 27369 96311
rect 27415 96265 27493 96311
rect 27539 96265 27617 96311
rect 27663 96265 27741 96311
rect 27787 96265 27865 96311
rect 27911 96265 27989 96311
rect 28035 96265 28113 96311
rect 28159 96265 28237 96311
rect 28283 96265 28361 96311
rect 28407 96265 28485 96311
rect 28531 96265 28609 96311
rect 28655 96265 28733 96311
rect 28779 96265 28857 96311
rect 28903 96265 28981 96311
rect 29027 96265 29105 96311
rect 29151 96265 29229 96311
rect 29275 96265 29353 96311
rect 29399 96265 29477 96311
rect 29523 96265 29601 96311
rect 29647 96265 29725 96311
rect 29771 96265 29849 96311
rect 29895 96265 29973 96311
rect 30019 96265 30097 96311
rect 30143 96265 30221 96311
rect 30267 96265 30345 96311
rect 30391 96265 30469 96311
rect 30515 96265 30593 96311
rect 30639 96265 30717 96311
rect 30763 96265 30841 96311
rect 30887 96265 30965 96311
rect 31011 96265 31089 96311
rect 31135 96265 31213 96311
rect 31259 96265 31337 96311
rect 31383 96265 31461 96311
rect 31507 96265 31585 96311
rect 31631 96265 31709 96311
rect 31755 96265 31833 96311
rect 31879 96265 31957 96311
rect 32003 96265 32081 96311
rect 32127 96265 32205 96311
rect 32251 96265 32329 96311
rect 32375 96265 32453 96311
rect 32499 96265 32577 96311
rect 32623 96265 32701 96311
rect 32747 96265 32825 96311
rect 32871 96265 32949 96311
rect 32995 96265 33073 96311
rect 33119 96265 33197 96311
rect 33243 96265 33321 96311
rect 33367 96265 33445 96311
rect 33491 96265 33569 96311
rect 33615 96265 33693 96311
rect 33739 96265 33817 96311
rect 33863 96265 33941 96311
rect 33987 96265 34065 96311
rect 34111 96265 34189 96311
rect 34235 96265 34313 96311
rect 34359 96265 34437 96311
rect 34483 96265 34561 96311
rect 34607 96265 34685 96311
rect 34731 96265 34809 96311
rect 34855 96265 34933 96311
rect 34979 96265 35057 96311
rect 35103 96265 35181 96311
rect 35227 96265 35305 96311
rect 35351 96265 35429 96311
rect 35475 96265 35553 96311
rect 35599 96265 35677 96311
rect 35723 96265 35801 96311
rect 35847 96265 35925 96311
rect 35971 96265 36049 96311
rect 36095 96265 36173 96311
rect 36219 96265 36297 96311
rect 36343 96265 36421 96311
rect 36467 96265 36545 96311
rect 36591 96265 36669 96311
rect 36715 96265 36793 96311
rect 36839 96265 36917 96311
rect 36963 96265 37041 96311
rect 37087 96265 37165 96311
rect 37211 96265 37289 96311
rect 37335 96265 37413 96311
rect 37459 96265 37537 96311
rect 37583 96265 37661 96311
rect 37707 96265 37785 96311
rect 37831 96265 37909 96311
rect 37955 96265 38033 96311
rect 38079 96265 38157 96311
rect 38203 96265 38281 96311
rect 38327 96265 38405 96311
rect 38451 96265 38529 96311
rect 38575 96265 38653 96311
rect 38699 96265 38777 96311
rect 38823 96265 38901 96311
rect 38947 96265 39025 96311
rect 39071 96265 39149 96311
rect 39195 96265 39273 96311
rect 39319 96265 39397 96311
rect 39443 96265 39521 96311
rect 39567 96265 39645 96311
rect 39691 96265 39769 96311
rect 39815 96265 39893 96311
rect 39939 96265 40017 96311
rect 40063 96265 40141 96311
rect 40187 96265 40265 96311
rect 40311 96265 40389 96311
rect 40435 96265 40513 96311
rect 40559 96265 40637 96311
rect 40683 96265 40761 96311
rect 40807 96265 40885 96311
rect 40931 96265 41009 96311
rect 41055 96265 41133 96311
rect 41179 96265 41257 96311
rect 41303 96265 41381 96311
rect 41427 96265 41505 96311
rect 41551 96265 41629 96311
rect 41675 96265 41753 96311
rect 41799 96265 41877 96311
rect 41923 96265 42001 96311
rect 42047 96265 42125 96311
rect 42171 96265 42249 96311
rect 42295 96265 42373 96311
rect 42419 96265 42497 96311
rect 42543 96265 42621 96311
rect 42667 96265 42745 96311
rect 42791 96265 42869 96311
rect 42915 96265 42993 96311
rect 43039 96265 43117 96311
rect 43163 96265 43241 96311
rect 43287 96265 43365 96311
rect 43411 96265 43489 96311
rect 43535 96265 43613 96311
rect 43659 96265 43737 96311
rect 43783 96265 43861 96311
rect 43907 96265 43985 96311
rect 44031 96265 44109 96311
rect 44155 96265 44233 96311
rect 44279 96265 44357 96311
rect 44403 96265 44481 96311
rect 44527 96265 44605 96311
rect 44651 96265 44729 96311
rect 44775 96265 44853 96311
rect 44899 96265 44977 96311
rect 45023 96265 45101 96311
rect 45147 96265 45225 96311
rect 45271 96265 45349 96311
rect 45395 96265 45473 96311
rect 45519 96265 45597 96311
rect 45643 96265 45721 96311
rect 45767 96265 45845 96311
rect 45891 96265 45969 96311
rect 46015 96265 46093 96311
rect 46139 96265 46217 96311
rect 46263 96265 46341 96311
rect 46387 96265 46465 96311
rect 46511 96265 46589 96311
rect 46635 96265 46713 96311
rect 46759 96265 46837 96311
rect 46883 96265 46961 96311
rect 47007 96265 47085 96311
rect 47131 96265 47209 96311
rect 47255 96265 47333 96311
rect 47379 96265 47457 96311
rect 47503 96265 47581 96311
rect 47627 96265 47705 96311
rect 47751 96265 47829 96311
rect 47875 96265 47953 96311
rect 47999 96265 48077 96311
rect 48123 96265 48201 96311
rect 48247 96265 48325 96311
rect 48371 96265 48449 96311
rect 48495 96265 48573 96311
rect 48619 96265 48697 96311
rect 48743 96265 48821 96311
rect 48867 96265 48945 96311
rect 48991 96265 49069 96311
rect 49115 96265 49193 96311
rect 49239 96265 49317 96311
rect 49363 96265 49441 96311
rect 49487 96265 49565 96311
rect 49611 96265 49689 96311
rect 49735 96265 49813 96311
rect 49859 96265 49937 96311
rect 49983 96265 50061 96311
rect 50107 96265 50185 96311
rect 50231 96265 50309 96311
rect 50355 96265 50433 96311
rect 50479 96265 50557 96311
rect 50603 96265 50681 96311
rect 50727 96265 50805 96311
rect 50851 96265 50929 96311
rect 50975 96265 51053 96311
rect 51099 96265 51177 96311
rect 51223 96265 51301 96311
rect 51347 96265 51425 96311
rect 51471 96265 51549 96311
rect 51595 96265 51673 96311
rect 51719 96265 51797 96311
rect 51843 96265 51921 96311
rect 51967 96265 52045 96311
rect 52091 96265 52169 96311
rect 52215 96265 52293 96311
rect 52339 96265 52417 96311
rect 52463 96265 52541 96311
rect 52587 96265 52665 96311
rect 52711 96265 52789 96311
rect 52835 96265 52913 96311
rect 52959 96265 53037 96311
rect 53083 96265 53161 96311
rect 53207 96265 53285 96311
rect 53331 96265 53409 96311
rect 53455 96265 53533 96311
rect 53579 96265 53657 96311
rect 53703 96265 53781 96311
rect 53827 96265 53905 96311
rect 53951 96265 54029 96311
rect 54075 96265 54153 96311
rect 54199 96265 54277 96311
rect 54323 96265 54401 96311
rect 54447 96265 54525 96311
rect 54571 96265 54649 96311
rect 54695 96265 54773 96311
rect 54819 96265 54897 96311
rect 54943 96265 55021 96311
rect 55067 96265 55145 96311
rect 55191 96265 55269 96311
rect 55315 96265 55393 96311
rect 55439 96265 55517 96311
rect 55563 96265 55641 96311
rect 55687 96265 55765 96311
rect 55811 96265 55889 96311
rect 55935 96265 56013 96311
rect 56059 96265 56137 96311
rect 56183 96265 56261 96311
rect 56307 96265 56385 96311
rect 56431 96265 56509 96311
rect 56555 96265 56633 96311
rect 56679 96265 56757 96311
rect 56803 96265 56881 96311
rect 56927 96265 57005 96311
rect 57051 96265 57129 96311
rect 57175 96265 57253 96311
rect 57299 96265 57377 96311
rect 57423 96265 57501 96311
rect 57547 96265 57625 96311
rect 57671 96265 57749 96311
rect 57795 96265 57873 96311
rect 57919 96265 57997 96311
rect 58043 96265 58121 96311
rect 58167 96265 58245 96311
rect 58291 96265 58369 96311
rect 58415 96265 58493 96311
rect 58539 96265 58617 96311
rect 58663 96265 58741 96311
rect 58787 96265 58865 96311
rect 58911 96265 58989 96311
rect 59035 96265 59113 96311
rect 59159 96265 59237 96311
rect 59283 96265 59361 96311
rect 59407 96265 59485 96311
rect 59531 96265 59609 96311
rect 59655 96265 59733 96311
rect 59779 96265 59857 96311
rect 59903 96265 59981 96311
rect 60027 96265 60105 96311
rect 60151 96265 60229 96311
rect 60275 96265 60353 96311
rect 60399 96265 60477 96311
rect 60523 96265 60601 96311
rect 60647 96265 60725 96311
rect 60771 96265 60849 96311
rect 60895 96265 60973 96311
rect 61019 96265 61097 96311
rect 61143 96265 61221 96311
rect 61267 96265 61345 96311
rect 61391 96265 61469 96311
rect 61515 96265 61593 96311
rect 61639 96265 61717 96311
rect 61763 96265 61841 96311
rect 61887 96265 61965 96311
rect 62011 96265 62089 96311
rect 62135 96265 62213 96311
rect 62259 96265 62337 96311
rect 62383 96265 62461 96311
rect 62507 96265 62585 96311
rect 62631 96265 62709 96311
rect 62755 96265 62833 96311
rect 62879 96265 62957 96311
rect 63003 96265 63081 96311
rect 63127 96265 63205 96311
rect 63251 96265 63329 96311
rect 63375 96265 63453 96311
rect 63499 96265 63577 96311
rect 63623 96265 63701 96311
rect 63747 96265 63825 96311
rect 63871 96265 63949 96311
rect 63995 96265 64073 96311
rect 64119 96265 64197 96311
rect 64243 96265 64321 96311
rect 64367 96265 64445 96311
rect 64491 96265 64569 96311
rect 64615 96265 64693 96311
rect 64739 96265 64817 96311
rect 64863 96265 64941 96311
rect 64987 96265 65065 96311
rect 65111 96265 65189 96311
rect 65235 96265 65313 96311
rect 65359 96265 65437 96311
rect 65483 96265 65561 96311
rect 65607 96265 65685 96311
rect 65731 96265 65809 96311
rect 65855 96265 65933 96311
rect 65979 96265 66057 96311
rect 66103 96265 66181 96311
rect 66227 96265 66305 96311
rect 66351 96265 66429 96311
rect 66475 96265 66553 96311
rect 66599 96265 66677 96311
rect 66723 96265 66801 96311
rect 66847 96265 66925 96311
rect 66971 96265 67049 96311
rect 67095 96265 67173 96311
rect 67219 96265 67297 96311
rect 67343 96265 67421 96311
rect 67467 96265 67545 96311
rect 67591 96265 67669 96311
rect 67715 96265 67793 96311
rect 67839 96265 67917 96311
rect 67963 96265 68041 96311
rect 68087 96265 68165 96311
rect 68211 96265 68289 96311
rect 68335 96265 68413 96311
rect 68459 96265 68537 96311
rect 68583 96265 68661 96311
rect 68707 96265 68785 96311
rect 68831 96265 68909 96311
rect 68955 96265 69033 96311
rect 69079 96265 69157 96311
rect 69203 96265 69281 96311
rect 69327 96265 69405 96311
rect 69451 96265 69529 96311
rect 69575 96265 69653 96311
rect 69699 96265 69777 96311
rect 69823 96265 69901 96311
rect 69947 96265 70025 96311
rect 70071 96265 70149 96311
rect 70195 96265 70273 96311
rect 70319 96265 70397 96311
rect 70443 96265 70521 96311
rect 70567 96265 70645 96311
rect 70691 96265 70769 96311
rect 70815 96265 70893 96311
rect 70939 96265 71017 96311
rect 71063 96265 71141 96311
rect 71187 96265 71265 96311
rect 71311 96265 71389 96311
rect 71435 96265 71513 96311
rect 71559 96265 71637 96311
rect 71683 96265 71761 96311
rect 71807 96265 71885 96311
rect 71931 96265 72009 96311
rect 72055 96265 72133 96311
rect 72179 96265 72257 96311
rect 72303 96265 72381 96311
rect 72427 96265 72505 96311
rect 72551 96265 72629 96311
rect 72675 96265 72753 96311
rect 72799 96265 72877 96311
rect 72923 96265 73001 96311
rect 73047 96265 73125 96311
rect 73171 96265 73249 96311
rect 73295 96265 73373 96311
rect 73419 96265 73497 96311
rect 73543 96265 73621 96311
rect 73667 96265 73745 96311
rect 73791 96265 73869 96311
rect 73915 96265 73993 96311
rect 74039 96265 74117 96311
rect 74163 96265 74241 96311
rect 74287 96265 74365 96311
rect 74411 96265 74489 96311
rect 74535 96265 74613 96311
rect 74659 96265 74737 96311
rect 74783 96265 74861 96311
rect 74907 96265 74985 96311
rect 75031 96265 75109 96311
rect 75155 96265 75233 96311
rect 75279 96265 75357 96311
rect 75403 96265 75481 96311
rect 75527 96265 75605 96311
rect 75651 96265 75729 96311
rect 75775 96265 75853 96311
rect 75899 96265 75977 96311
rect 76023 96265 76101 96311
rect 76147 96265 76225 96311
rect 76271 96265 76349 96311
rect 76395 96265 76473 96311
rect 76519 96265 76597 96311
rect 76643 96265 76721 96311
rect 76767 96265 76845 96311
rect 76891 96265 76969 96311
rect 77015 96265 77093 96311
rect 77139 96265 77217 96311
rect 77263 96265 77341 96311
rect 77387 96265 77465 96311
rect 77511 96265 77589 96311
rect 77635 96265 77713 96311
rect 77759 96265 77837 96311
rect 77883 96265 77961 96311
rect 78007 96265 78085 96311
rect 78131 96265 78209 96311
rect 78255 96265 78333 96311
rect 78379 96265 78457 96311
rect 78503 96265 78581 96311
rect 78627 96265 78705 96311
rect 78751 96265 78829 96311
rect 78875 96265 78953 96311
rect 78999 96265 79077 96311
rect 79123 96265 79201 96311
rect 79247 96265 79325 96311
rect 79371 96265 79449 96311
rect 79495 96265 79573 96311
rect 79619 96265 79697 96311
rect 79743 96265 79821 96311
rect 79867 96265 79945 96311
rect 79991 96265 80069 96311
rect 80115 96265 80193 96311
rect 80239 96265 80317 96311
rect 80363 96265 80441 96311
rect 80487 96265 80565 96311
rect 80611 96265 80689 96311
rect 80735 96265 80813 96311
rect 80859 96265 80937 96311
rect 80983 96265 81061 96311
rect 81107 96265 81185 96311
rect 81231 96265 81309 96311
rect 81355 96265 81433 96311
rect 81479 96265 81557 96311
rect 81603 96265 81681 96311
rect 81727 96265 81805 96311
rect 81851 96265 81929 96311
rect 81975 96265 82053 96311
rect 82099 96265 82177 96311
rect 82223 96265 82301 96311
rect 82347 96265 82425 96311
rect 82471 96265 82549 96311
rect 82595 96265 82673 96311
rect 82719 96265 82797 96311
rect 82843 96265 82921 96311
rect 82967 96265 83045 96311
rect 83091 96265 83169 96311
rect 83215 96265 83293 96311
rect 83339 96265 83417 96311
rect 83463 96265 83541 96311
rect 83587 96265 83665 96311
rect 83711 96265 83789 96311
rect 83835 96265 83913 96311
rect 83959 96265 84037 96311
rect 84083 96265 84161 96311
rect 84207 96265 84285 96311
rect 84331 96265 84409 96311
rect 84455 96265 84533 96311
rect 84579 96265 84657 96311
rect 84703 96265 84781 96311
rect 84827 96265 84905 96311
rect 84951 96265 85029 96311
rect 85075 96265 85153 96311
rect 85199 96265 85277 96311
rect 85323 96265 85401 96311
rect 85447 96265 85525 96311
rect 85571 96265 85649 96311
rect 85695 96265 85706 96311
rect 0 96254 85706 96265
rect 0 96163 1000 96254
rect 0 1117 89 96163
rect 435 1117 1000 96163
rect 0 1026 1000 1117
rect 27105 96163 27473 96174
rect 27105 1117 27116 96163
rect 27462 1117 27473 96163
rect 57013 96163 57381 96174
rect 27529 96142 28397 96153
rect 27529 35996 27540 96142
rect 28386 35996 28397 96142
rect 27529 35985 28397 35996
rect 56089 96142 56957 96153
rect 56089 35996 56100 96142
rect 56946 35996 56957 96142
rect 56089 35985 56957 35996
rect 27529 34620 56897 34631
rect 27529 34174 27540 34620
rect 56886 34174 56897 34620
rect 27529 34163 56897 34174
rect 27105 1106 27473 1117
rect 57013 1117 57024 96163
rect 57370 1117 57381 96163
rect 57013 1106 57381 1117
rect 85440 96163 85808 96174
rect 85440 1117 85451 96163
rect 85797 1117 85808 96163
rect 85440 1106 85808 1117
rect 0 1015 85706 1026
rect 0 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85706 1015
rect 0 891 85706 969
rect 0 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85706 891
rect 0 767 85706 845
rect 0 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85706 767
rect 0 643 85706 721
rect 0 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85706 643
rect 0 586 85706 597
rect 0 403 1000 586
<< metal2 >>
rect 424 403 1424 96149
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_0
timestamp 1755724134
transform -1 0 85672 0 1 96288
box 0 0 1 1
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_1
timestamp 1755724134
transform -1 0 85672 0 1 620
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_0
timestamp 1755724134
transform 1 0 85474 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_1
timestamp 1755724134
transform 1 0 27139 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_2
timestamp 1755724134
transform 1 0 57047 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_3
timestamp 1755724134
transform 1 0 112 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_0
timestamp 1755724134
transform 1 0 56123 0 1 36019
box 0 0 1 1
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_1
timestamp 1755724134
transform 1 0 27563 0 1 36019
box 0 0 1 1
use M1_PSUB4310591302046_512x8m81  M1_PSUB4310591302046_512x8m81_0
timestamp 1755724134
transform 1 0 27563 0 1 34197
box 0 0 1 1
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 448 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2641664
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2640354
string path 4.620 11.160 4.620 0.000 
<< end >>
