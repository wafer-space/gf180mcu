magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 4118 1094
<< pwell >>
rect -86 -86 4118 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 179 836 297
rect 940 179 1060 297
rect 1164 179 1284 297
rect 1332 179 1452 297
rect 1624 215 1744 333
rect 1808 215 1928 333
rect 2032 215 2152 333
rect 2256 215 2376 333
rect 2872 215 2992 333
rect 3056 215 3176 333
rect 3324 183 3444 333
rect 3692 69 3812 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 736 593 836 793
rect 960 593 1060 793
rect 1164 593 1264 793
rect 1332 593 1432 793
rect 1624 593 1724 793
rect 1828 593 1928 793
rect 2256 573 2356 773
rect 2524 573 2624 773
rect 2872 593 2972 793
rect 3076 593 3176 793
rect 3316 573 3416 793
rect 3712 573 3812 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 1544 297 1624 333
rect 468 175 556 274
rect 628 238 716 297
rect 628 192 641 238
rect 687 192 716 238
rect 628 179 716 192
rect 836 284 940 297
rect 836 238 865 284
rect 911 238 940 284
rect 836 179 940 238
rect 1060 284 1164 297
rect 1060 238 1089 284
rect 1135 238 1164 284
rect 1060 179 1164 238
rect 1284 179 1332 297
rect 1452 238 1624 297
rect 1452 192 1481 238
rect 1527 215 1624 238
rect 1744 215 1808 333
rect 1928 320 2032 333
rect 1928 274 1957 320
rect 2003 274 2032 320
rect 1928 215 2032 274
rect 2152 274 2256 333
rect 2152 228 2181 274
rect 2227 228 2256 274
rect 2152 215 2256 228
rect 2376 320 2464 333
rect 2376 274 2405 320
rect 2451 274 2464 320
rect 2376 215 2464 274
rect 1527 192 1540 215
rect 1452 179 1540 192
rect 2784 309 2872 333
rect 2784 263 2797 309
rect 2843 263 2872 309
rect 2784 215 2872 263
rect 2992 215 3056 333
rect 3176 242 3324 333
rect 3176 215 3249 242
rect 3236 196 3249 215
rect 3295 196 3324 242
rect 3236 183 3324 196
rect 3444 320 3532 333
rect 3444 274 3473 320
rect 3519 274 3532 320
rect 3444 183 3532 274
rect 3604 222 3692 333
rect 3604 82 3617 222
rect 3663 82 3692 222
rect 3604 69 3692 82
rect 3812 320 3900 333
rect 3812 180 3841 320
rect 3887 180 3900 320
rect 3812 69 3900 180
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 1492 943 1564 956
rect 1492 803 1505 943
rect 1551 803 1564 943
rect 1492 793 1564 803
rect 1988 858 2060 871
rect 1988 812 2001 858
rect 2047 812 2060 858
rect 1988 793 2060 812
rect 448 586 477 726
rect 523 586 536 726
rect 648 780 736 793
rect 648 640 661 780
rect 707 640 736 780
rect 648 593 736 640
rect 836 746 960 793
rect 836 606 865 746
rect 911 606 960 746
rect 836 593 960 606
rect 1060 746 1164 793
rect 1060 606 1089 746
rect 1135 606 1164 746
rect 1060 593 1164 606
rect 1264 593 1332 793
rect 1432 593 1624 793
rect 1724 652 1828 793
rect 1724 606 1753 652
rect 1799 606 1828 652
rect 1724 593 1828 606
rect 1928 593 2060 793
rect 3624 926 3712 939
rect 2784 780 2872 793
rect 2168 652 2256 773
rect 2168 606 2181 652
rect 2227 606 2256 652
rect 448 573 536 586
rect 2168 573 2256 606
rect 2356 726 2524 773
rect 2356 586 2385 726
rect 2431 586 2524 726
rect 2356 573 2524 586
rect 2624 726 2712 773
rect 2624 586 2653 726
rect 2699 586 2712 726
rect 2784 640 2797 780
rect 2843 640 2872 780
rect 2784 593 2872 640
rect 2972 746 3076 793
rect 2972 606 3001 746
rect 3047 606 3076 746
rect 2972 593 3076 606
rect 3176 780 3316 793
rect 3176 734 3205 780
rect 3251 734 3316 780
rect 3176 593 3316 734
rect 2624 573 2712 586
rect 3236 573 3316 593
rect 3416 632 3504 793
rect 3416 586 3445 632
rect 3491 586 3504 632
rect 3416 573 3504 586
rect 3624 786 3637 926
rect 3683 786 3712 926
rect 3624 573 3712 786
rect 3812 726 3900 939
rect 3812 586 3841 726
rect 3887 586 3900 726
rect 3812 573 3900 586
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 192 687 238
rect 865 238 911 284
rect 1089 238 1135 284
rect 1481 192 1527 238
rect 1957 274 2003 320
rect 2181 228 2227 274
rect 2405 274 2451 320
rect 2797 263 2843 309
rect 3249 196 3295 242
rect 3473 274 3519 320
rect 3617 82 3663 222
rect 3841 180 3887 320
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 1505 803 1551 943
rect 2001 812 2047 858
rect 477 586 523 726
rect 661 640 707 780
rect 865 606 911 746
rect 1089 606 1135 746
rect 1753 606 1799 652
rect 2181 606 2227 652
rect 2385 586 2431 726
rect 2653 586 2699 726
rect 2797 640 2843 780
rect 3001 606 3047 746
rect 3205 734 3251 780
rect 3445 586 3491 632
rect 3637 786 3683 926
rect 3841 586 3887 726
<< polysilicon >>
rect 348 933 1264 973
rect 144 849 244 893
rect 348 849 448 933
rect 960 872 1060 885
rect 736 793 836 837
rect 960 826 973 872
rect 1019 826 1060 872
rect 960 793 1060 826
rect 1164 872 1264 933
rect 1164 826 1205 872
rect 1251 826 1264 872
rect 1164 793 1264 826
rect 1332 793 1432 837
rect 1828 931 2972 971
rect 3712 939 3812 983
rect 1624 793 1724 837
rect 1828 793 1928 931
rect 2256 852 2356 865
rect 2256 806 2269 852
rect 2315 806 2356 852
rect 2256 773 2356 806
rect 2524 773 2624 817
rect 2872 793 2972 931
rect 3076 793 3176 837
rect 3316 793 3416 837
rect 144 512 244 573
rect 144 466 157 512
rect 203 466 244 512
rect 144 377 244 466
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 736 400 836 593
rect 960 504 1060 593
rect 1164 549 1264 593
rect 1332 560 1432 593
rect 1332 514 1373 560
rect 1419 514 1432 560
rect 960 464 1147 504
rect 407 366 468 377
rect 348 333 468 366
rect 736 354 749 400
rect 795 354 836 400
rect 1107 397 1147 464
rect 1107 376 1284 397
rect 1107 357 1225 376
rect 736 341 836 354
rect 716 297 836 341
rect 940 297 1060 341
rect 1164 330 1225 357
rect 1271 330 1284 376
rect 1164 297 1284 330
rect 1332 341 1432 514
rect 1624 468 1724 593
rect 1624 422 1637 468
rect 1683 422 1724 468
rect 1624 377 1724 422
rect 1828 377 1928 593
rect 2256 377 2356 573
rect 1332 297 1452 341
rect 1624 333 1744 377
rect 1808 333 1928 377
rect 2032 333 2152 377
rect 2256 333 2376 377
rect 124 131 244 175
rect 348 87 468 175
rect 716 135 836 179
rect 940 87 1060 179
rect 1164 135 1284 179
rect 1332 135 1452 179
rect 1624 171 1744 215
rect 1808 171 1928 215
rect 2032 182 2152 215
rect 2032 136 2045 182
rect 2091 136 2152 182
rect 2256 171 2376 215
rect 348 47 1060 87
rect 2032 123 2152 136
rect 2524 123 2624 573
rect 2872 423 2972 593
rect 2872 377 2885 423
rect 2931 377 2972 423
rect 3076 560 3176 593
rect 3076 514 3117 560
rect 3163 514 3176 560
rect 3076 377 3176 514
rect 3316 412 3416 573
rect 3316 393 3337 412
rect 2872 333 2992 377
rect 3056 333 3176 377
rect 3324 366 3337 393
rect 3383 393 3416 412
rect 3712 535 3812 573
rect 3712 489 3725 535
rect 3771 489 3812 535
rect 3383 366 3444 393
rect 3712 377 3812 489
rect 3324 333 3444 366
rect 3692 333 3812 377
rect 2872 171 2992 215
rect 3056 171 3176 215
rect 3324 139 3444 183
rect 2032 83 2624 123
rect 3692 25 3812 69
<< polycontact >>
rect 973 826 1019 872
rect 1205 826 1251 872
rect 2269 806 2315 852
rect 157 466 203 512
rect 361 366 407 412
rect 1373 514 1419 560
rect 749 354 795 400
rect 1225 330 1271 376
rect 1637 422 1683 468
rect 2045 136 2091 182
rect 2885 377 2931 423
rect 3117 514 3163 560
rect 3337 366 3383 412
rect 3725 489 3771 535
<< metal1 >>
rect 0 943 4032 1098
rect 0 918 1505 943
rect 273 836 319 918
rect 69 739 115 750
rect 661 780 707 918
rect 273 685 319 696
rect 477 726 523 737
rect 115 599 407 634
rect 69 588 407 599
rect 142 512 306 542
rect 142 466 157 512
rect 203 466 306 512
rect 361 412 407 588
rect 49 366 361 401
rect 49 355 407 366
rect 661 629 707 640
rect 753 826 973 872
rect 1019 826 1030 872
rect 1194 826 1205 872
rect 1251 826 1262 872
rect 477 583 523 586
rect 753 583 799 826
rect 477 537 799 583
rect 865 746 911 757
rect 49 320 95 355
rect 49 263 95 274
rect 477 320 543 537
rect 590 400 806 430
rect 590 354 749 400
rect 795 354 806 400
rect 477 274 497 320
rect 477 263 543 274
rect 865 284 911 606
rect 273 234 319 245
rect 273 90 319 188
rect 641 238 687 249
rect 865 227 911 238
rect 1089 746 1135 757
rect 1194 746 1262 826
rect 1551 926 4032 943
rect 1551 918 3637 926
rect 1505 792 1551 803
rect 2001 858 2047 918
rect 2001 801 2047 812
rect 2269 852 2315 863
rect 2269 755 2315 806
rect 1579 746 2315 755
rect 1194 709 2315 746
rect 2797 780 2843 918
rect 2385 726 2431 737
rect 1194 700 1607 709
rect 1089 468 1135 606
rect 1753 652 2227 663
rect 1799 606 2181 652
rect 1753 595 2227 606
rect 1753 560 2003 595
rect 1362 514 1373 560
rect 1419 514 2003 560
rect 1089 422 1637 468
rect 1683 422 1694 468
rect 1089 284 1135 422
rect 1214 330 1225 376
rect 1271 330 1619 376
rect 1089 227 1135 238
rect 1481 238 1527 249
rect 641 90 687 192
rect 1481 90 1527 192
rect 1573 182 1619 330
rect 1957 320 2003 514
rect 2385 423 2431 586
rect 2653 726 2699 737
rect 3205 780 3251 918
rect 2797 629 2843 640
rect 3001 746 3047 757
rect 2653 583 2699 586
rect 3683 918 4032 926
rect 3637 775 3683 786
rect 3205 723 3251 734
rect 3838 726 3890 737
rect 3001 583 3047 606
rect 2653 537 3047 583
rect 3117 632 3491 643
rect 3117 586 3445 632
rect 3117 560 3491 586
rect 2653 526 2699 537
rect 1957 263 2003 274
rect 2181 377 2431 423
rect 2502 480 2699 526
rect 3163 546 3491 560
rect 3838 586 3841 726
rect 3887 586 3890 726
rect 3163 535 3771 546
rect 3163 514 3725 535
rect 3117 503 3725 514
rect 3473 489 3725 503
rect 2181 274 2227 377
rect 2502 331 2548 480
rect 3473 478 3771 489
rect 2594 423 2931 434
rect 2594 377 2885 423
rect 2594 366 2931 377
rect 2977 366 3337 412
rect 3383 366 3394 412
rect 2405 320 2548 331
rect 2451 309 2843 320
rect 2451 274 2797 309
rect 2405 263 2797 274
rect 2405 252 2843 263
rect 2181 206 2227 228
rect 2977 206 3023 366
rect 3473 320 3519 478
rect 3473 263 3519 274
rect 3838 320 3890 586
rect 1573 136 2045 182
rect 2091 136 2102 182
rect 2181 160 3023 206
rect 3249 242 3295 253
rect 3249 90 3295 196
rect 3617 222 3663 233
rect 0 82 3617 90
rect 3838 180 3841 320
rect 3887 180 3890 320
rect 3838 169 3890 180
rect 3663 82 4032 90
rect 0 -90 4032 82
<< labels >>
flabel metal1 s 142 466 306 542 0 FreeSans 200 0 0 0 CLK
port 3 nsew clock input
flabel metal1 s 590 354 806 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3838 169 3890 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2594 366 2931 434 0 FreeSans 200 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 918 4032 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3249 249 3295 253 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3637 801 3683 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3205 801 3251 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 801 2843 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2001 801 2047 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1505 801 1551 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 801 707 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 801 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3637 792 3683 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3205 792 3251 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 792 2843 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1505 792 1551 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 792 707 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 792 319 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3637 775 3683 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3205 775 3251 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 775 2843 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 775 707 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3205 723 3251 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 723 2843 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 723 707 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 723 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 685 2843 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 685 707 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2797 629 2843 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 629 707 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3249 245 3295 249 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1481 245 1527 249 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 245 687 249 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3249 233 3295 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1481 233 1527 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3617 90 3663 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3249 90 3295 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1481 90 1527 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4032 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 1008
string GDS_END 673602
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 664556
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
