magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 377 4902 870
rect -86 352 1889 377
rect 4588 352 4902 377
<< pwell >>
rect -86 -86 4902 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 2060 93 2180 257
rect 2284 93 2404 257
rect 2508 93 2628 257
rect 2732 93 2852 257
rect 2956 93 3076 257
rect 3180 93 3300 257
rect 3404 93 3524 257
rect 3628 93 3748 257
rect 3852 93 3972 257
rect 4076 93 4196 257
rect 4300 93 4420 257
rect 4568 68 4688 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 572 497 672 716
rect 816 497 916 716
rect 1020 497 1120 716
rect 1264 497 1364 716
rect 1468 497 1568 716
rect 1712 497 1812 716
rect 2080 529 2180 716
rect 2284 529 2384 716
rect 2528 529 2628 716
rect 2732 529 2832 716
rect 2976 497 3076 716
rect 3200 497 3300 716
rect 3404 497 3504 716
rect 3648 497 3748 716
rect 3852 497 3952 716
rect 4096 497 4196 716
rect 4300 497 4400 716
rect 4568 497 4668 716
<< mvndiff >>
rect 36 127 124 232
rect 36 81 49 127
rect 95 81 124 127
rect 36 68 124 81
rect 244 219 348 232
rect 244 173 273 219
rect 319 173 348 219
rect 244 68 348 173
rect 468 127 572 232
rect 468 81 497 127
rect 543 81 572 127
rect 468 68 572 81
rect 692 219 796 232
rect 692 173 721 219
rect 767 173 796 219
rect 692 68 796 173
rect 916 127 1020 232
rect 916 81 945 127
rect 991 81 1020 127
rect 916 68 1020 81
rect 1140 219 1244 232
rect 1140 173 1169 219
rect 1215 173 1244 219
rect 1140 68 1244 173
rect 1364 127 1468 232
rect 1364 81 1393 127
rect 1439 81 1468 127
rect 1364 68 1468 81
rect 1588 219 1692 232
rect 1588 173 1617 219
rect 1663 173 1692 219
rect 1588 68 1692 173
rect 1812 127 1900 232
rect 1812 81 1841 127
rect 1887 81 1900 127
rect 1972 152 2060 257
rect 1972 106 1985 152
rect 2031 106 2060 152
rect 1972 93 2060 106
rect 2180 244 2284 257
rect 2180 198 2209 244
rect 2255 198 2284 244
rect 2180 93 2284 198
rect 2404 152 2508 257
rect 2404 106 2433 152
rect 2479 106 2508 152
rect 2404 93 2508 106
rect 2628 244 2732 257
rect 2628 198 2657 244
rect 2703 198 2732 244
rect 2628 93 2732 198
rect 2852 152 2956 257
rect 2852 106 2881 152
rect 2927 106 2956 152
rect 2852 93 2956 106
rect 3076 244 3180 257
rect 3076 198 3105 244
rect 3151 198 3180 244
rect 3076 93 3180 198
rect 3300 152 3404 257
rect 3300 106 3329 152
rect 3375 106 3404 152
rect 3300 93 3404 106
rect 3524 244 3628 257
rect 3524 198 3553 244
rect 3599 198 3628 244
rect 3524 93 3628 198
rect 3748 152 3852 257
rect 3748 106 3777 152
rect 3823 106 3852 152
rect 3748 93 3852 106
rect 3972 244 4076 257
rect 3972 198 4001 244
rect 4047 198 4076 244
rect 3972 93 4076 198
rect 4196 152 4300 257
rect 4196 106 4225 152
rect 4271 106 4300 152
rect 4196 93 4300 106
rect 4420 244 4508 257
rect 4420 198 4449 244
rect 4495 232 4508 244
rect 4495 198 4568 232
rect 4420 93 4568 198
rect 1812 68 1900 81
rect 4488 68 4568 93
rect 4688 152 4776 232
rect 4688 106 4717 152
rect 4763 106 4776 152
rect 4688 68 4776 106
<< mvpdiff >>
rect 56 611 144 716
rect 56 565 69 611
rect 115 565 144 611
rect 56 497 144 565
rect 244 497 368 716
rect 468 664 572 716
rect 468 618 497 664
rect 543 618 572 664
rect 468 497 572 618
rect 672 497 816 716
rect 916 611 1020 716
rect 916 565 945 611
rect 991 565 1020 611
rect 916 497 1020 565
rect 1120 497 1264 716
rect 1364 664 1468 716
rect 1364 618 1393 664
rect 1439 618 1468 664
rect 1364 497 1468 618
rect 1568 497 1712 716
rect 1812 611 2080 716
rect 1812 565 1841 611
rect 1887 565 2005 611
rect 2051 565 2080 611
rect 1812 529 2080 565
rect 2180 664 2284 716
rect 2180 618 2209 664
rect 2255 618 2284 664
rect 2180 529 2284 618
rect 2384 611 2528 716
rect 2384 565 2433 611
rect 2479 565 2528 611
rect 2384 529 2528 565
rect 2628 664 2732 716
rect 2628 618 2657 664
rect 2703 618 2732 664
rect 2628 529 2732 618
rect 2832 611 2976 716
rect 2832 565 2881 611
rect 2927 565 2976 611
rect 2832 529 2976 565
rect 1812 497 1912 529
rect 2896 497 2976 529
rect 3076 497 3200 716
rect 3300 703 3404 716
rect 3300 657 3329 703
rect 3375 657 3404 703
rect 3300 497 3404 657
rect 3504 497 3648 716
rect 3748 662 3852 716
rect 3748 616 3777 662
rect 3823 616 3852 662
rect 3748 497 3852 616
rect 3952 497 4096 716
rect 4196 703 4300 716
rect 4196 657 4225 703
rect 4271 657 4300 703
rect 4196 497 4300 657
rect 4400 497 4568 716
rect 4668 611 4756 716
rect 4668 565 4697 611
rect 4743 565 4756 611
rect 4668 497 4756 565
<< mvndiffc >>
rect 49 81 95 127
rect 273 173 319 219
rect 497 81 543 127
rect 721 173 767 219
rect 945 81 991 127
rect 1169 173 1215 219
rect 1393 81 1439 127
rect 1617 173 1663 219
rect 1841 81 1887 127
rect 1985 106 2031 152
rect 2209 198 2255 244
rect 2433 106 2479 152
rect 2657 198 2703 244
rect 2881 106 2927 152
rect 3105 198 3151 244
rect 3329 106 3375 152
rect 3553 198 3599 244
rect 3777 106 3823 152
rect 4001 198 4047 244
rect 4225 106 4271 152
rect 4449 198 4495 244
rect 4717 106 4763 152
<< mvpdiffc >>
rect 69 565 115 611
rect 497 618 543 664
rect 945 565 991 611
rect 1393 618 1439 664
rect 1841 565 1887 611
rect 2005 565 2051 611
rect 2209 618 2255 664
rect 2433 565 2479 611
rect 2657 618 2703 664
rect 2881 565 2927 611
rect 3329 657 3375 703
rect 3777 616 3823 662
rect 4225 657 4271 703
rect 4697 565 4743 611
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 1020 716 1120 760
rect 1264 716 1364 760
rect 1468 716 1568 760
rect 1712 716 1812 760
rect 2080 716 2180 760
rect 2284 716 2384 760
rect 2528 716 2628 760
rect 2732 716 2832 760
rect 2976 716 3076 760
rect 3200 716 3300 760
rect 3404 716 3504 760
rect 3648 716 3748 760
rect 3852 716 3952 760
rect 4096 716 4196 760
rect 4300 716 4400 760
rect 4568 716 4668 760
rect 144 415 244 497
rect 144 402 171 415
rect 124 369 171 402
rect 217 369 244 415
rect 368 415 468 497
rect 368 402 395 415
rect 124 232 244 369
rect 348 369 395 402
rect 441 394 468 415
rect 572 415 672 497
rect 572 394 599 415
rect 441 369 599 394
rect 645 402 672 415
rect 816 402 916 497
rect 645 369 692 402
rect 348 348 692 369
rect 348 232 468 348
rect 572 232 692 348
rect 796 394 916 402
rect 1020 402 1120 497
rect 1264 415 1364 497
rect 1264 402 1291 415
rect 1020 394 1140 402
rect 796 348 1140 394
rect 796 314 916 348
rect 796 268 833 314
rect 879 268 916 314
rect 796 232 916 268
rect 1020 314 1140 348
rect 1020 268 1057 314
rect 1103 268 1140 314
rect 1020 232 1140 268
rect 1244 369 1291 402
rect 1337 394 1364 415
rect 1468 415 1568 497
rect 1468 394 1485 415
rect 1337 369 1485 394
rect 1531 402 1568 415
rect 1712 415 1812 497
rect 1712 402 1739 415
rect 1531 369 1588 402
rect 1244 348 1588 369
rect 1244 232 1364 348
rect 1468 232 1588 348
rect 1692 369 1739 402
rect 1785 369 1812 415
rect 2080 415 2180 529
rect 2080 402 2107 415
rect 1692 232 1812 369
rect 2060 369 2107 402
rect 2153 402 2180 415
rect 2284 415 2384 529
rect 2284 402 2311 415
rect 2153 369 2311 402
rect 2357 402 2384 415
rect 2528 415 2628 529
rect 2528 402 2555 415
rect 2357 369 2555 402
rect 2601 402 2628 415
rect 2732 415 2832 529
rect 2732 402 2759 415
rect 2601 369 2759 402
rect 2805 402 2832 415
rect 2976 402 3076 497
rect 3200 415 3300 497
rect 3200 402 3227 415
rect 2805 369 2852 402
rect 2060 348 2852 369
rect 2060 257 2180 348
rect 2284 257 2404 348
rect 2508 257 2628 348
rect 2732 257 2852 348
rect 2956 394 3076 402
rect 2956 348 3003 394
rect 3049 348 3076 394
rect 2956 257 3076 348
rect 3180 369 3227 402
rect 3273 394 3300 415
rect 3404 415 3504 497
rect 3404 394 3431 415
rect 3273 369 3431 394
rect 3477 402 3504 415
rect 3648 428 3748 497
rect 3648 402 3675 428
rect 3477 369 3524 402
rect 3180 348 3524 369
rect 3180 257 3300 348
rect 3404 257 3524 348
rect 3628 382 3675 402
rect 3721 394 3748 428
rect 3852 428 3952 497
rect 3852 394 3879 428
rect 3721 382 3879 394
rect 3925 402 3952 428
rect 4096 402 4196 497
rect 3925 382 3972 402
rect 3628 348 3972 382
rect 3628 257 3748 348
rect 3852 257 3972 348
rect 4076 394 4196 402
rect 4300 402 4400 497
rect 4568 418 4668 497
rect 4300 394 4420 402
rect 4076 348 4420 394
rect 4076 336 4196 348
rect 4076 290 4113 336
rect 4159 290 4196 336
rect 4076 257 4196 290
rect 4300 336 4420 348
rect 4300 290 4319 336
rect 4365 290 4420 336
rect 4300 257 4420 290
rect 4568 372 4595 418
rect 4641 402 4668 418
rect 4641 372 4688 402
rect 4568 232 4688 372
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 2060 24 2180 93
rect 2284 24 2404 93
rect 2508 24 2628 93
rect 2732 24 2852 93
rect 2956 24 3076 93
rect 3180 24 3300 93
rect 3404 24 3524 93
rect 3628 24 3748 93
rect 3852 24 3972 93
rect 4076 24 4196 93
rect 4300 24 4420 93
rect 4568 24 4688 68
<< polycontact >>
rect 171 369 217 415
rect 395 369 441 415
rect 599 369 645 415
rect 833 268 879 314
rect 1057 268 1103 314
rect 1291 369 1337 415
rect 1485 369 1531 415
rect 1739 369 1785 415
rect 2107 369 2153 415
rect 2311 369 2357 415
rect 2555 369 2601 415
rect 2759 369 2805 415
rect 3003 348 3049 394
rect 3227 369 3273 415
rect 3431 369 3477 415
rect 3675 382 3721 428
rect 3879 382 3925 428
rect 4113 290 4159 336
rect 4319 290 4365 336
rect 4595 372 4641 418
<< metal1 >>
rect 0 724 4816 844
rect 486 664 554 724
rect 69 611 115 622
rect 486 618 497 664
rect 543 618 554 664
rect 1382 664 1450 724
rect 69 536 115 565
rect 945 611 991 622
rect 1382 618 1393 664
rect 1439 618 1450 664
rect 2198 664 2266 724
rect 945 536 991 565
rect 1841 611 1887 622
rect 1841 536 1887 565
rect 2005 611 2051 622
rect 2198 618 2209 664
rect 2255 618 2266 664
rect 2646 664 2714 724
rect 2005 536 2051 565
rect 2433 611 2479 622
rect 2646 618 2657 664
rect 2703 618 2714 664
rect 3318 703 3386 724
rect 3318 657 3329 703
rect 3375 657 3386 703
rect 4214 703 4282 724
rect 3447 616 3777 662
rect 3823 616 4147 662
rect 4214 657 4225 703
rect 4271 657 4282 703
rect 3447 611 4147 616
rect 2433 536 2479 565
rect 2870 565 2881 611
rect 2927 582 4697 611
rect 2927 565 3493 582
rect 4101 565 4697 582
rect 4743 565 4756 611
rect 2870 536 2938 565
rect 69 472 2938 536
rect 3594 519 4022 536
rect 124 415 318 424
rect 124 369 171 415
rect 217 369 318 415
rect 124 360 318 369
rect 368 415 1542 424
rect 368 369 395 415
rect 441 369 599 415
rect 645 369 1291 415
rect 1337 369 1485 415
rect 1531 369 1542 415
rect 368 360 1542 369
rect 1588 415 1894 424
rect 1588 369 1739 415
rect 1785 369 1894 415
rect 270 314 318 360
rect 1588 354 1894 369
rect 2023 415 2832 424
rect 2023 369 2107 415
rect 2153 369 2311 415
rect 2357 369 2555 415
rect 2601 369 2759 415
rect 2805 369 2832 415
rect 2023 360 2832 369
rect 1588 314 1634 354
rect 270 268 833 314
rect 879 268 1057 314
rect 1103 268 1634 314
rect 2881 244 2938 472
rect 3003 473 4022 519
rect 3003 394 3049 473
rect 3664 428 3732 473
rect 3143 415 3585 424
rect 3143 369 3227 415
rect 3273 369 3431 415
rect 3477 369 3585 415
rect 3664 382 3675 428
rect 3721 382 3732 428
rect 3868 428 4022 473
rect 3868 382 3879 428
rect 3925 418 4684 428
rect 3925 382 4595 418
rect 3143 360 3585 369
rect 3003 320 3049 348
rect 3535 336 3585 360
rect 4477 372 4595 382
rect 4641 372 4684 418
rect 4477 358 4684 372
rect 3535 290 4113 336
rect 4159 290 4319 336
rect 4365 290 4376 336
rect 1757 219 2209 244
rect 244 173 273 219
rect 319 173 721 219
rect 767 173 1169 219
rect 1215 173 1617 219
rect 1663 198 2209 219
rect 2255 198 2657 244
rect 2703 198 2714 244
rect 2881 198 3105 244
rect 3151 198 3553 244
rect 3599 198 4001 244
rect 4047 198 4449 244
rect 4495 198 4506 244
rect 4612 224 4684 358
rect 1663 173 1807 198
rect 38 81 49 127
rect 95 81 106 127
rect 38 60 106 81
rect 485 81 497 127
rect 543 81 554 127
rect 485 60 554 81
rect 933 81 945 127
rect 991 81 1002 127
rect 933 60 1002 81
rect 1381 81 1393 127
rect 1439 81 1450 127
rect 1381 60 1450 81
rect 1829 81 1841 127
rect 1887 81 1898 127
rect 1972 106 1985 152
rect 2031 106 2433 152
rect 2479 106 2881 152
rect 2927 106 3329 152
rect 3375 106 3777 152
rect 3823 106 4225 152
rect 4271 106 4717 152
rect 4763 106 4776 152
rect 1829 60 1898 81
rect 0 -60 4816 60
<< labels >>
flabel metal1 s 3594 519 4022 536 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1588 360 1894 424 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 368 360 1542 424 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel metal1 s 2023 360 2832 424 0 FreeSans 400 0 0 0 C
port 5 nsew default input
flabel metal1 s 0 724 4816 844 0 FreeSans 400 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 1829 60 1898 127 0 FreeSans 400 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 3447 622 4147 662 0 FreeSans 400 0 0 0 ZN
port 6 nsew default output
flabel metal1 s 3143 360 3585 424 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 8 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 3003 473 4022 519 1 A1
port 1 nsew default input
rlabel metal1 s 3868 428 4022 473 1 A1
port 1 nsew default input
rlabel metal1 s 3664 428 3732 473 1 A1
port 1 nsew default input
rlabel metal1 s 3003 428 3049 473 1 A1
port 1 nsew default input
rlabel metal1 s 3868 382 4684 428 1 A1
port 1 nsew default input
rlabel metal1 s 3664 382 3732 428 1 A1
port 1 nsew default input
rlabel metal1 s 3003 382 3049 428 1 A1
port 1 nsew default input
rlabel metal1 s 4477 358 4684 382 1 A1
port 1 nsew default input
rlabel metal1 s 3003 358 3049 382 1 A1
port 1 nsew default input
rlabel metal1 s 4612 320 4684 358 1 A1
port 1 nsew default input
rlabel metal1 s 3003 320 3049 358 1 A1
port 1 nsew default input
rlabel metal1 s 4612 224 4684 320 1 A1
port 1 nsew default input
rlabel metal1 s 3535 336 3585 360 1 A2
port 2 nsew default input
rlabel metal1 s 3535 290 4376 336 1 A2
port 2 nsew default input
rlabel metal1 s 124 360 318 424 1 B1
port 3 nsew default input
rlabel metal1 s 1588 354 1894 360 1 B1
port 3 nsew default input
rlabel metal1 s 270 354 318 360 1 B1
port 3 nsew default input
rlabel metal1 s 1588 314 1634 354 1 B1
port 3 nsew default input
rlabel metal1 s 270 314 318 354 1 B1
port 3 nsew default input
rlabel metal1 s 270 268 1634 314 1 B1
port 3 nsew default input
rlabel metal1 s 3447 611 4147 622 1 ZN
port 6 nsew default output
rlabel metal1 s 2433 611 2479 622 1 ZN
port 6 nsew default output
rlabel metal1 s 2005 611 2051 622 1 ZN
port 6 nsew default output
rlabel metal1 s 1841 611 1887 622 1 ZN
port 6 nsew default output
rlabel metal1 s 945 611 991 622 1 ZN
port 6 nsew default output
rlabel metal1 s 69 611 115 622 1 ZN
port 6 nsew default output
rlabel metal1 s 2870 582 4756 611 1 ZN
port 6 nsew default output
rlabel metal1 s 2433 582 2479 611 1 ZN
port 6 nsew default output
rlabel metal1 s 2005 582 2051 611 1 ZN
port 6 nsew default output
rlabel metal1 s 1841 582 1887 611 1 ZN
port 6 nsew default output
rlabel metal1 s 945 582 991 611 1 ZN
port 6 nsew default output
rlabel metal1 s 69 582 115 611 1 ZN
port 6 nsew default output
rlabel metal1 s 4101 565 4756 582 1 ZN
port 6 nsew default output
rlabel metal1 s 2870 565 3493 582 1 ZN
port 6 nsew default output
rlabel metal1 s 2433 565 2479 582 1 ZN
port 6 nsew default output
rlabel metal1 s 2005 565 2051 582 1 ZN
port 6 nsew default output
rlabel metal1 s 1841 565 1887 582 1 ZN
port 6 nsew default output
rlabel metal1 s 945 565 991 582 1 ZN
port 6 nsew default output
rlabel metal1 s 69 565 115 582 1 ZN
port 6 nsew default output
rlabel metal1 s 2870 536 2938 565 1 ZN
port 6 nsew default output
rlabel metal1 s 2433 536 2479 565 1 ZN
port 6 nsew default output
rlabel metal1 s 2005 536 2051 565 1 ZN
port 6 nsew default output
rlabel metal1 s 1841 536 1887 565 1 ZN
port 6 nsew default output
rlabel metal1 s 945 536 991 565 1 ZN
port 6 nsew default output
rlabel metal1 s 69 536 115 565 1 ZN
port 6 nsew default output
rlabel metal1 s 69 472 2938 536 1 ZN
port 6 nsew default output
rlabel metal1 s 2881 244 2938 472 1 ZN
port 6 nsew default output
rlabel metal1 s 2881 198 4506 244 1 ZN
port 6 nsew default output
rlabel metal1 s 4214 657 4282 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3318 657 3386 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2646 657 2714 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2198 657 2266 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1382 657 1450 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 486 657 554 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2646 618 2714 657 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2198 618 2266 657 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1382 618 1450 657 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 486 618 554 657 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1381 60 1450 127 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 933 60 1002 127 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 485 60 554 127 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 127 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4816 60 1 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 784
string GDS_END 123072
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 114708
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
