magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< mvnmos >>
rect 124 156 244 296
rect 348 156 468 296
rect 572 156 692 296
rect 796 156 916 296
rect 964 156 1084 296
rect 1188 156 1308 296
rect 1556 161 1676 301
rect 1780 161 1900 301
rect 2236 161 2356 321
rect 2460 161 2580 321
rect 2684 161 2804 321
rect 3116 133 3236 333
rect 3340 133 3460 333
<< mvpmos >>
rect 362 576 462 852
rect 510 576 610 852
rect 680 576 780 852
rect 884 576 984 852
rect 1032 576 1132 852
rect 1236 576 1336 852
rect 1596 573 1696 849
rect 1800 573 1900 849
rect 2276 573 2376 909
rect 2480 573 2580 909
rect 2628 573 2728 909
rect 3126 573 3226 939
rect 3330 573 3430 939
<< mvndiff >>
rect 36 220 124 296
rect 36 174 49 220
rect 95 174 124 220
rect 36 156 124 174
rect 244 220 348 296
rect 244 174 273 220
rect 319 174 348 220
rect 244 156 348 174
rect 468 220 572 296
rect 468 174 497 220
rect 543 174 572 220
rect 468 156 572 174
rect 692 220 796 296
rect 692 174 721 220
rect 767 174 796 220
rect 692 156 796 174
rect 916 156 964 296
rect 1084 220 1188 296
rect 1084 174 1113 220
rect 1159 174 1188 220
rect 1084 156 1188 174
rect 1308 220 1396 296
rect 1308 174 1337 220
rect 1383 174 1396 220
rect 1308 156 1396 174
rect 1468 220 1556 301
rect 1468 174 1481 220
rect 1527 174 1556 220
rect 1468 161 1556 174
rect 1676 220 1780 301
rect 1676 174 1705 220
rect 1751 174 1780 220
rect 1676 161 1780 174
rect 1900 220 1988 301
rect 1900 174 1929 220
rect 1975 174 1988 220
rect 1900 161 1988 174
rect 2148 308 2236 321
rect 2148 262 2161 308
rect 2207 262 2236 308
rect 2148 161 2236 262
rect 2356 220 2460 321
rect 2356 174 2385 220
rect 2431 174 2460 220
rect 2356 161 2460 174
rect 2580 308 2684 321
rect 2580 262 2609 308
rect 2655 262 2684 308
rect 2580 161 2684 262
rect 2804 220 2892 321
rect 2804 174 2833 220
rect 2879 174 2892 220
rect 2804 161 2892 174
rect 3028 314 3116 333
rect 3028 174 3041 314
rect 3087 174 3116 314
rect 3028 133 3116 174
rect 3236 314 3340 333
rect 3236 174 3265 314
rect 3311 174 3340 314
rect 3236 133 3340 174
rect 3460 314 3548 333
rect 3460 174 3489 314
rect 3535 174 3548 314
rect 3460 133 3548 174
<< mvpdiff >>
rect 274 831 362 852
rect 274 691 287 831
rect 333 691 362 831
rect 274 576 362 691
rect 462 576 510 852
rect 610 576 680 852
rect 780 831 884 852
rect 780 691 809 831
rect 855 691 884 831
rect 780 576 884 691
rect 984 576 1032 852
rect 1132 831 1236 852
rect 1132 691 1161 831
rect 1207 691 1236 831
rect 1132 576 1236 691
rect 1336 769 1424 852
rect 1336 629 1365 769
rect 1411 629 1424 769
rect 1336 576 1424 629
rect 1508 769 1596 849
rect 1508 629 1521 769
rect 1567 629 1596 769
rect 1508 573 1596 629
rect 1696 831 1800 849
rect 1696 691 1725 831
rect 1771 691 1800 831
rect 1696 573 1800 691
rect 1900 831 1988 849
rect 1900 691 1929 831
rect 1975 691 1988 831
rect 1900 573 1988 691
rect 2188 733 2276 909
rect 2188 593 2201 733
rect 2247 593 2276 733
rect 2188 573 2276 593
rect 2376 831 2480 909
rect 2376 691 2405 831
rect 2451 691 2480 831
rect 2376 573 2480 691
rect 2580 573 2628 909
rect 2728 831 2816 909
rect 2728 691 2757 831
rect 2803 691 2816 831
rect 2728 573 2816 691
rect 3038 831 3126 939
rect 3038 691 3051 831
rect 3097 691 3126 831
rect 3038 573 3126 691
rect 3226 831 3330 939
rect 3226 691 3255 831
rect 3301 691 3330 831
rect 3226 573 3330 691
rect 3430 831 3518 939
rect 3430 691 3459 831
rect 3505 691 3518 831
rect 3430 573 3518 691
<< mvndiffc >>
rect 49 174 95 220
rect 273 174 319 220
rect 497 174 543 220
rect 721 174 767 220
rect 1113 174 1159 220
rect 1337 174 1383 220
rect 1481 174 1527 220
rect 1705 174 1751 220
rect 1929 174 1975 220
rect 2161 262 2207 308
rect 2385 174 2431 220
rect 2609 262 2655 308
rect 2833 174 2879 220
rect 3041 174 3087 314
rect 3265 174 3311 314
rect 3489 174 3535 314
<< mvpdiffc >>
rect 287 691 333 831
rect 809 691 855 831
rect 1161 691 1207 831
rect 1365 629 1411 769
rect 1521 629 1567 769
rect 1725 691 1771 831
rect 1929 691 1975 831
rect 2201 593 2247 733
rect 2405 691 2451 831
rect 2757 691 2803 831
rect 3051 691 3097 831
rect 3255 691 3301 831
rect 3459 691 3505 831
<< polysilicon >>
rect 1032 944 1900 984
rect 362 852 462 896
rect 510 852 610 896
rect 680 852 780 896
rect 884 852 984 896
rect 1032 852 1132 944
rect 1236 852 1336 896
rect 1596 849 1696 893
rect 1800 849 1900 944
rect 2276 909 2376 953
rect 2480 909 2580 953
rect 2628 909 2728 953
rect 3126 939 3226 983
rect 3330 939 3430 983
rect 362 532 462 576
rect 510 532 610 576
rect 680 532 780 576
rect 362 509 402 532
rect 335 471 402 509
rect 335 447 375 471
rect 510 447 550 532
rect 740 516 780 532
rect 884 542 984 576
rect 740 476 836 516
rect 884 496 898 542
rect 944 496 984 542
rect 884 483 984 496
rect 1032 532 1132 576
rect 1236 532 1336 576
rect 124 434 375 447
rect 124 388 148 434
rect 194 407 375 434
rect 444 434 550 447
rect 444 407 478 434
rect 194 388 244 407
rect 124 296 244 388
rect 428 388 478 407
rect 524 419 550 434
rect 524 388 539 419
rect 428 375 539 388
rect 652 415 748 428
rect 428 340 468 375
rect 652 369 689 415
rect 735 369 748 415
rect 652 356 748 369
rect 652 340 692 356
rect 348 296 468 340
rect 572 296 692 340
rect 796 340 836 476
rect 1032 340 1084 532
rect 1236 340 1308 532
rect 1596 434 1696 573
rect 1596 388 1623 434
rect 1669 388 1696 434
rect 1596 377 1696 388
rect 1800 434 1900 573
rect 2276 531 2376 573
rect 2276 485 2289 531
rect 2335 529 2376 531
rect 2480 540 2580 573
rect 2335 485 2356 529
rect 1800 388 1813 434
rect 1859 388 1900 434
rect 1596 345 1676 377
rect 1800 345 1900 388
rect 796 296 916 340
rect 964 296 1084 340
rect 1188 296 1308 340
rect 1556 301 1676 345
rect 1780 301 1900 345
rect 2048 434 2120 447
rect 2048 388 2061 434
rect 2107 388 2120 434
rect 2048 375 2120 388
rect 124 112 244 156
rect 348 112 468 156
rect 572 112 692 156
rect 796 64 916 156
rect 964 112 1084 156
rect 1188 64 1308 156
rect 1556 117 1676 161
rect 1780 117 1900 161
rect 2048 64 2088 375
rect 2276 365 2356 485
rect 2480 494 2493 540
rect 2539 494 2580 540
rect 2628 529 2728 573
rect 2480 365 2580 494
rect 2236 321 2356 365
rect 2460 321 2580 365
rect 2684 365 2728 529
rect 3126 465 3226 573
rect 3330 465 3430 573
rect 3126 434 3430 465
rect 3126 388 3139 434
rect 3185 393 3430 434
rect 3185 388 3236 393
rect 3126 377 3236 388
rect 2684 321 2804 365
rect 3116 333 3236 377
rect 3340 377 3430 393
rect 3340 333 3460 377
rect 796 24 2088 64
rect 2236 69 2356 161
rect 2460 117 2580 161
rect 2684 69 2804 161
rect 3116 89 3236 133
rect 3340 89 3460 133
rect 2236 29 2804 69
<< polycontact >>
rect 898 496 944 542
rect 148 388 194 434
rect 478 388 524 434
rect 689 369 735 415
rect 1623 388 1669 434
rect 2289 485 2335 531
rect 1813 388 1859 434
rect 2061 388 2107 434
rect 2493 494 2539 540
rect 3139 388 3185 434
<< metal1 >>
rect 0 918 3584 1098
rect 287 831 333 918
rect 287 680 333 691
rect 809 831 855 842
rect 809 634 855 691
rect 1161 831 1207 918
rect 1161 680 1207 691
rect 1253 826 1669 872
rect 1253 634 1299 826
rect 809 613 1299 634
rect 586 588 1299 613
rect 1365 769 1411 780
rect 586 567 848 588
rect 142 434 194 542
rect 142 388 148 434
rect 142 354 194 388
rect 478 434 530 542
rect 524 388 530 434
rect 478 354 530 388
rect 586 323 632 567
rect 887 496 898 542
rect 944 496 955 542
rect 887 415 955 496
rect 1365 415 1411 629
rect 678 369 689 415
rect 735 369 1411 415
rect 213 308 459 312
rect 49 266 459 308
rect 586 277 767 323
rect 49 262 232 266
rect 49 220 95 262
rect 413 231 459 266
rect 413 220 543 231
rect 49 163 95 174
rect 262 174 273 220
rect 319 174 330 220
rect 262 90 330 174
rect 413 174 497 220
rect 413 163 543 174
rect 721 220 767 277
rect 721 163 767 174
rect 1113 220 1159 231
rect 1113 90 1159 174
rect 1337 220 1411 369
rect 1383 174 1411 220
rect 1337 163 1411 174
rect 1481 769 1567 780
rect 1481 629 1521 769
rect 1481 331 1567 629
rect 1623 434 1669 826
rect 1725 831 1771 918
rect 1725 680 1771 691
rect 1929 831 2359 842
rect 1975 796 2359 831
rect 1623 377 1669 388
rect 1715 388 1813 434
rect 1859 388 1870 434
rect 1715 331 1761 388
rect 1481 285 1761 331
rect 1481 220 1527 285
rect 1481 163 1527 174
rect 1705 220 1751 231
rect 1705 90 1751 174
rect 1929 220 1975 691
rect 2201 733 2247 744
rect 2061 593 2201 628
rect 2061 582 2247 593
rect 2313 634 2359 796
rect 2405 831 2451 918
rect 2405 680 2451 691
rect 2757 831 2803 842
rect 2313 588 2539 634
rect 2061 434 2107 582
rect 2061 308 2107 388
rect 2270 531 2335 542
rect 2270 485 2289 531
rect 2270 354 2335 485
rect 2493 540 2539 588
rect 2493 483 2539 494
rect 2757 434 2803 691
rect 3051 831 3097 918
rect 3051 680 3097 691
rect 3255 831 3330 842
rect 3301 691 3330 831
rect 2757 388 3139 434
rect 3185 388 3196 434
rect 2757 312 2803 388
rect 2598 308 2803 312
rect 2061 262 2161 308
rect 2207 262 2218 308
rect 2598 262 2609 308
rect 2655 266 2803 308
rect 3041 314 3087 325
rect 2655 262 2666 266
rect 1929 163 1975 174
rect 2385 220 2431 231
rect 2385 90 2431 174
rect 2833 220 2879 231
rect 2833 90 2879 174
rect 3041 90 3087 174
rect 3255 314 3330 691
rect 3459 831 3505 918
rect 3459 680 3505 691
rect 3255 174 3265 314
rect 3311 174 3330 314
rect 3255 163 3330 174
rect 3489 314 3535 325
rect 3489 90 3535 174
rect 0 -90 3584 90
<< labels >>
flabel metal1 s 2270 354 2335 542 0 FreeSans 200 0 0 0 CLKN
port 1 nsew clock input
flabel metal1 s 478 354 530 542 0 FreeSans 200 0 0 0 E
port 2 nsew default input
flabel metal1 s 3255 163 3330 842 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 918 3584 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3489 231 3535 325 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3459 680 3505 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3051 680 3097 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2405 680 2451 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1725 680 1771 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1161 680 1207 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 287 680 333 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3041 231 3087 325 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3489 220 3535 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3041 220 3087 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2833 220 2879 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2385 220 2431 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1705 220 1751 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1113 220 1159 231 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3489 90 3535 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3041 90 3087 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2833 90 2879 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2385 90 2431 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1705 90 1751 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1113 90 1159 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 220 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3584 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string GDS_END 835924
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 827488
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
