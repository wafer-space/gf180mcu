magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 534 870
<< pwell >>
rect -86 -86 534 352
<< mvnmos >>
rect 124 68 244 232
<< mvpmos >>
rect 144 472 244 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 244 192 332 232
rect 244 146 273 192
rect 319 146 332 192
rect 244 68 332 146
<< mvpdiff >>
rect 56 665 144 716
rect 56 525 69 665
rect 115 525 144 665
rect 56 472 144 525
rect 244 665 332 716
rect 244 525 273 665
rect 319 525 332 665
rect 244 472 332 525
<< mvndiffc >>
rect 49 146 95 192
rect 273 146 319 192
<< mvpdiffc >>
rect 69 525 115 665
rect 273 525 319 665
<< polysilicon >>
rect 144 716 244 760
rect 144 423 244 472
rect 144 386 157 423
rect 124 283 157 386
rect 203 283 244 423
rect 124 232 244 283
rect 124 24 244 68
<< polycontact >>
rect 157 283 203 423
<< metal1 >>
rect 0 724 448 844
rect 69 665 115 724
rect 69 506 115 525
rect 253 665 319 678
rect 253 525 273 665
rect 142 423 207 440
rect 142 283 157 423
rect 203 283 207 423
rect 142 240 207 283
rect 49 192 95 232
rect 49 60 95 146
rect 253 192 319 525
rect 253 146 273 192
rect 253 106 319 146
rect 0 -60 448 60
<< labels >>
flabel metal1 s 49 60 95 232 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 253 106 319 678 0 FreeSans 400 0 0 0 ZN
port 2 nsew default output
flabel metal1 s 142 240 207 440 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 448 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 69 506 115 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -60 448 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string GDS_END 476332
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 474136
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
