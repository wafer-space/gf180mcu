magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 1878 870
<< pwell >>
rect -86 -86 1878 352
<< metal1 >>
rect 0 724 1792 844
rect 253 632 299 724
rect 661 632 707 724
rect 869 472 1534 556
rect 124 364 806 424
rect 330 206 418 318
rect 869 230 944 472
rect 990 360 1676 424
rect 990 280 1047 360
rect 1138 242 1676 314
rect 49 60 95 181
rect 188 122 418 206
rect 464 220 944 230
rect 464 174 1031 220
rect 464 143 511 174
rect 985 128 1330 174
rect 854 60 922 128
rect 1681 60 1727 181
rect 0 -60 1792 60
<< obsm1 >>
rect 38 552 106 676
rect 446 552 514 676
rect 759 626 1738 673
rect 759 552 805 626
rect 38 506 805 552
rect 1670 495 1738 626
<< labels >>
rlabel metal1 s 1138 242 1676 314 6 A1
port 1 nsew default input
rlabel metal1 s 990 280 1047 360 6 A2
port 2 nsew default input
rlabel metal1 s 990 360 1676 424 6 A2
port 2 nsew default input
rlabel metal1 s 188 122 418 206 6 B1
port 3 nsew default input
rlabel metal1 s 330 206 418 318 6 B1
port 3 nsew default input
rlabel metal1 s 124 364 806 424 6 B2
port 4 nsew default input
rlabel metal1 s 985 128 1330 174 6 ZN
port 5 nsew default output
rlabel metal1 s 464 143 511 174 6 ZN
port 5 nsew default output
rlabel metal1 s 464 174 1031 220 6 ZN
port 5 nsew default output
rlabel metal1 s 464 220 944 230 6 ZN
port 5 nsew default output
rlabel metal1 s 869 230 944 472 6 ZN
port 5 nsew default output
rlabel metal1 s 869 472 1534 556 6 ZN
port 5 nsew default output
rlabel metal1 s 661 632 707 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 632 299 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 724 1792 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel nwell s -86 352 1878 870 6 VNW
port 7 nsew power bidirectional
rlabel pwell s -86 -86 1878 352 6 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 0 -60 1792 60 8 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1681 60 1727 181 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 854 60 922 128 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 181 6 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1269246
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1264704
<< end >>
