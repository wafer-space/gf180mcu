magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 6470 1094
<< pwell >>
rect -86 -86 6470 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 978 68 1098 332
rect 1202 68 1322 332
rect 1426 68 1546 332
rect 1650 68 1770 332
rect 1874 68 1994 332
rect 2098 68 2218 332
rect 2322 68 2442 332
rect 2546 68 2666 332
rect 2770 68 2890 332
rect 2994 68 3114 332
rect 3218 68 3338 332
rect 3442 68 3562 332
rect 3666 68 3786 332
rect 3890 68 4010 332
rect 4114 68 4234 332
rect 4338 68 4458 332
rect 4562 68 4682 332
rect 4786 68 4906 332
rect 5010 68 5130 332
rect 5234 68 5354 332
rect 5458 68 5578 332
rect 5682 68 5802 332
rect 5906 68 6026 332
rect 6130 68 6250 332
<< mvpmos >>
rect 172 573 272 933
rect 376 573 476 933
rect 660 573 760 933
rect 1058 573 1158 933
rect 1262 573 1362 933
rect 1466 573 1566 933
rect 1670 573 1770 933
rect 1874 573 1974 933
rect 2138 573 2238 933
rect 2342 573 2442 933
rect 2582 580 2682 940
rect 2786 580 2886 940
rect 2990 580 3090 940
rect 3194 580 3294 940
rect 3398 580 3498 940
rect 3602 580 3702 940
rect 3806 580 3906 940
rect 4010 580 4110 940
rect 4214 580 4314 940
rect 4418 580 4518 940
rect 4622 580 4722 940
rect 4826 580 4926 940
rect 5030 580 5130 940
rect 5234 580 5334 940
rect 5438 580 5538 940
rect 5642 580 5742 940
rect 5846 580 5946 940
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 69 124 274
rect 244 128 348 333
rect 244 82 273 128
rect 319 82 348 128
rect 244 69 348 82
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 320 780 333
rect 692 274 721 320
rect 767 274 780 320
rect 692 69 780 274
rect 852 125 978 332
rect 852 79 865 125
rect 911 79 978 125
rect 852 68 978 79
rect 1098 272 1202 332
rect 1098 226 1127 272
rect 1173 226 1202 272
rect 1098 68 1202 226
rect 1322 127 1426 332
rect 1322 81 1351 127
rect 1397 81 1426 127
rect 1322 68 1426 81
rect 1546 319 1650 332
rect 1546 179 1575 319
rect 1621 179 1650 319
rect 1546 68 1650 179
rect 1770 127 1874 332
rect 1770 81 1799 127
rect 1845 81 1874 127
rect 1770 68 1874 81
rect 1994 319 2098 332
rect 1994 179 2023 319
rect 2069 179 2098 319
rect 1994 68 2098 179
rect 2218 127 2322 332
rect 2218 81 2247 127
rect 2293 81 2322 127
rect 2218 68 2322 81
rect 2442 319 2546 332
rect 2442 179 2471 319
rect 2517 179 2546 319
rect 2442 68 2546 179
rect 2666 127 2770 332
rect 2666 81 2695 127
rect 2741 81 2770 127
rect 2666 68 2770 81
rect 2890 272 2994 332
rect 2890 226 2919 272
rect 2965 226 2994 272
rect 2890 68 2994 226
rect 3114 127 3218 332
rect 3114 81 3143 127
rect 3189 81 3218 127
rect 3114 68 3218 81
rect 3338 319 3442 332
rect 3338 179 3367 319
rect 3413 179 3442 319
rect 3338 68 3442 179
rect 3562 127 3666 332
rect 3562 81 3591 127
rect 3637 81 3666 127
rect 3562 68 3666 81
rect 3786 319 3890 332
rect 3786 179 3815 319
rect 3861 179 3890 319
rect 3786 68 3890 179
rect 4010 127 4114 332
rect 4010 81 4039 127
rect 4085 81 4114 127
rect 4010 68 4114 81
rect 4234 319 4338 332
rect 4234 179 4263 319
rect 4309 179 4338 319
rect 4234 68 4338 179
rect 4458 127 4562 332
rect 4458 81 4487 127
rect 4533 81 4562 127
rect 4458 68 4562 81
rect 4682 319 4786 332
rect 4682 179 4711 319
rect 4757 179 4786 319
rect 4682 68 4786 179
rect 4906 127 5010 332
rect 4906 81 4935 127
rect 4981 81 5010 127
rect 4906 68 5010 81
rect 5130 319 5234 332
rect 5130 179 5159 319
rect 5205 179 5234 319
rect 5130 68 5234 179
rect 5354 127 5458 332
rect 5354 81 5383 127
rect 5429 81 5458 127
rect 5354 68 5458 81
rect 5578 319 5682 332
rect 5578 179 5607 319
rect 5653 179 5682 319
rect 5578 68 5682 179
rect 5802 127 5906 332
rect 5802 81 5831 127
rect 5877 81 5906 127
rect 5802 68 5906 81
rect 6026 272 6130 332
rect 6026 226 6055 272
rect 6101 226 6130 272
rect 6026 68 6130 226
rect 6250 221 6338 332
rect 6250 81 6279 221
rect 6325 81 6338 221
rect 6250 68 6338 81
rect 852 66 918 68
<< mvpdiff >>
rect 2502 933 2582 940
rect 84 739 172 933
rect 84 599 97 739
rect 143 599 172 739
rect 84 573 172 599
rect 272 920 376 933
rect 272 780 301 920
rect 347 780 376 920
rect 272 573 376 780
rect 476 771 660 933
rect 476 725 585 771
rect 631 725 660 771
rect 476 573 660 725
rect 760 632 848 933
rect 760 586 789 632
rect 835 586 848 632
rect 760 573 848 586
rect 970 920 1058 933
rect 970 874 983 920
rect 1029 874 1058 920
rect 970 573 1058 874
rect 1158 817 1262 933
rect 1158 677 1187 817
rect 1233 677 1262 817
rect 1158 573 1262 677
rect 1362 920 1466 933
rect 1362 874 1391 920
rect 1437 874 1466 920
rect 1362 573 1466 874
rect 1566 817 1670 933
rect 1566 677 1595 817
rect 1641 677 1670 817
rect 1566 573 1670 677
rect 1770 920 1874 933
rect 1770 874 1799 920
rect 1845 874 1874 920
rect 1770 573 1874 874
rect 1974 817 2138 933
rect 1974 677 2003 817
rect 2049 677 2138 817
rect 1974 573 2138 677
rect 2238 920 2342 933
rect 2238 874 2267 920
rect 2313 874 2342 920
rect 2238 573 2342 874
rect 2442 770 2582 933
rect 2442 724 2471 770
rect 2517 724 2582 770
rect 2442 580 2582 724
rect 2682 927 2786 940
rect 2682 881 2711 927
rect 2757 881 2786 927
rect 2682 580 2786 881
rect 2886 778 2990 940
rect 2886 732 2915 778
rect 2961 732 2990 778
rect 2886 580 2990 732
rect 3090 927 3194 940
rect 3090 881 3119 927
rect 3165 881 3194 927
rect 3090 580 3194 881
rect 3294 824 3398 940
rect 3294 684 3323 824
rect 3369 684 3398 824
rect 3294 580 3398 684
rect 3498 927 3602 940
rect 3498 881 3527 927
rect 3573 881 3602 927
rect 3498 580 3602 881
rect 3702 824 3806 940
rect 3702 684 3731 824
rect 3777 684 3806 824
rect 3702 580 3806 684
rect 3906 927 4010 940
rect 3906 881 3935 927
rect 3981 881 4010 927
rect 3906 580 4010 881
rect 4110 824 4214 940
rect 4110 684 4139 824
rect 4185 684 4214 824
rect 4110 580 4214 684
rect 4314 927 4418 940
rect 4314 881 4343 927
rect 4389 881 4418 927
rect 4314 580 4418 881
rect 4518 824 4622 940
rect 4518 684 4547 824
rect 4593 684 4622 824
rect 4518 580 4622 684
rect 4722 927 4826 940
rect 4722 881 4751 927
rect 4797 881 4826 927
rect 4722 580 4826 881
rect 4926 824 5030 940
rect 4926 684 4955 824
rect 5001 684 5030 824
rect 4926 580 5030 684
rect 5130 927 5234 940
rect 5130 881 5159 927
rect 5205 881 5234 927
rect 5130 580 5234 881
rect 5334 824 5438 940
rect 5334 684 5363 824
rect 5409 684 5438 824
rect 5334 580 5438 684
rect 5538 927 5642 940
rect 5538 881 5567 927
rect 5613 881 5642 927
rect 5538 580 5642 881
rect 5742 824 5846 940
rect 5742 684 5771 824
rect 5817 684 5846 824
rect 5742 580 5846 684
rect 5946 927 6034 940
rect 5946 787 5975 927
rect 6021 787 6034 927
rect 5946 580 6034 787
rect 2442 573 2522 580
<< mvndiffc >>
rect 49 274 95 320
rect 273 82 319 128
rect 497 147 543 287
rect 721 274 767 320
rect 865 79 911 125
rect 1127 226 1173 272
rect 1351 81 1397 127
rect 1575 179 1621 319
rect 1799 81 1845 127
rect 2023 179 2069 319
rect 2247 81 2293 127
rect 2471 179 2517 319
rect 2695 81 2741 127
rect 2919 226 2965 272
rect 3143 81 3189 127
rect 3367 179 3413 319
rect 3591 81 3637 127
rect 3815 179 3861 319
rect 4039 81 4085 127
rect 4263 179 4309 319
rect 4487 81 4533 127
rect 4711 179 4757 319
rect 4935 81 4981 127
rect 5159 179 5205 319
rect 5383 81 5429 127
rect 5607 179 5653 319
rect 5831 81 5877 127
rect 6055 226 6101 272
rect 6279 81 6325 221
<< mvpdiffc >>
rect 97 599 143 739
rect 301 780 347 920
rect 585 725 631 771
rect 789 586 835 632
rect 983 874 1029 920
rect 1187 677 1233 817
rect 1391 874 1437 920
rect 1595 677 1641 817
rect 1799 874 1845 920
rect 2003 677 2049 817
rect 2267 874 2313 920
rect 2471 724 2517 770
rect 2711 881 2757 927
rect 2915 732 2961 778
rect 3119 881 3165 927
rect 3323 684 3369 824
rect 3527 881 3573 927
rect 3731 684 3777 824
rect 3935 881 3981 927
rect 4139 684 4185 824
rect 4343 881 4389 927
rect 4547 684 4593 824
rect 4751 881 4797 927
rect 4955 684 5001 824
rect 5159 881 5205 927
rect 5363 684 5409 824
rect 5567 881 5613 927
rect 5771 684 5817 824
rect 5975 787 6021 927
<< polysilicon >>
rect 172 933 272 977
rect 376 933 476 977
rect 660 933 760 977
rect 1058 933 1158 977
rect 1262 933 1362 977
rect 1466 933 1566 977
rect 1670 933 1770 977
rect 1874 933 1974 977
rect 2138 933 2238 977
rect 2342 933 2442 977
rect 2582 940 2682 984
rect 2786 940 2886 984
rect 2990 940 3090 984
rect 3194 940 3294 984
rect 3398 940 3498 984
rect 3602 940 3702 984
rect 3806 940 3906 984
rect 4010 940 4110 984
rect 4214 940 4314 984
rect 4418 940 4518 984
rect 4622 940 4722 984
rect 4826 940 4926 984
rect 5030 940 5130 984
rect 5234 940 5334 984
rect 5438 940 5538 984
rect 5642 940 5742 984
rect 5846 940 5946 984
rect 172 523 272 573
rect 172 477 185 523
rect 231 513 272 523
rect 376 513 476 573
rect 660 540 760 573
rect 231 477 612 513
rect 660 494 673 540
rect 719 494 760 540
rect 660 481 760 494
rect 1058 509 1158 573
rect 172 473 612 477
rect 172 377 244 473
rect 124 333 244 377
rect 348 412 468 425
rect 348 366 361 412
rect 407 366 468 412
rect 348 333 468 366
rect 572 377 612 473
rect 1058 463 1085 509
rect 1131 473 1158 509
rect 1262 509 1362 573
rect 1262 473 1287 509
rect 1131 463 1287 473
rect 1333 473 1362 509
rect 1466 509 1566 573
rect 1466 473 1492 509
rect 1333 463 1492 473
rect 1538 473 1566 509
rect 1670 509 1770 573
rect 1670 473 1695 509
rect 1538 463 1695 473
rect 1741 473 1770 509
rect 1874 509 1974 573
rect 1874 473 1901 509
rect 1741 463 1901 473
rect 1947 473 1974 509
rect 2138 509 2238 573
rect 2138 473 2165 509
rect 1947 463 2165 473
rect 2211 473 2238 509
rect 2342 509 2442 573
rect 2342 473 2369 509
rect 2211 463 2369 473
rect 2415 473 2442 509
rect 2582 473 2682 580
rect 2786 540 2886 580
rect 2786 494 2816 540
rect 2862 520 2886 540
rect 2990 540 3090 580
rect 2990 520 3019 540
rect 2862 494 3019 520
rect 3065 520 3090 540
rect 3194 540 3294 580
rect 3194 520 3223 540
rect 3065 494 3223 520
rect 3269 520 3294 540
rect 3398 540 3498 580
rect 3398 520 3427 540
rect 3269 494 3427 520
rect 3473 520 3498 540
rect 3602 540 3702 580
rect 3602 520 3629 540
rect 3473 494 3629 520
rect 3675 520 3702 540
rect 3806 540 3906 580
rect 3806 520 3833 540
rect 3675 494 3833 520
rect 3879 520 3906 540
rect 4010 540 4110 580
rect 4010 520 4038 540
rect 3879 494 4038 520
rect 4084 520 4110 540
rect 4214 540 4314 580
rect 4214 520 4241 540
rect 4084 494 4241 520
rect 4287 520 4314 540
rect 4418 540 4518 580
rect 4418 520 4447 540
rect 4287 494 4447 520
rect 4493 520 4518 540
rect 4622 540 4722 580
rect 4622 520 4651 540
rect 4493 494 4651 520
rect 4697 520 4722 540
rect 4826 540 4926 580
rect 4826 520 4854 540
rect 4697 494 4854 520
rect 4900 520 4926 540
rect 5030 540 5130 580
rect 5030 520 5058 540
rect 4900 494 5058 520
rect 5104 520 5130 540
rect 5234 540 5334 580
rect 5234 520 5260 540
rect 5104 494 5260 520
rect 5306 520 5334 540
rect 5438 540 5538 580
rect 5438 520 5467 540
rect 5306 494 5467 520
rect 5513 520 5538 540
rect 5642 520 5742 580
rect 5846 520 5946 580
rect 5513 494 5946 520
rect 2786 480 5946 494
rect 2415 463 2682 473
rect 1058 433 2682 463
rect 572 333 692 377
rect 1058 376 1098 433
rect 978 332 1098 376
rect 1202 332 1322 433
rect 1426 332 1546 433
rect 1650 332 1770 433
rect 1874 332 1994 433
rect 2098 332 2218 433
rect 2322 332 2442 433
rect 2546 332 2666 433
rect 2770 419 6250 432
rect 2770 373 2783 419
rect 2829 392 3032 419
rect 2829 373 2890 392
rect 2770 332 2890 373
rect 2994 373 3032 392
rect 3078 392 3255 419
rect 3078 373 3114 392
rect 2994 332 3114 373
rect 3218 373 3255 392
rect 3301 392 3478 419
rect 3301 373 3338 392
rect 3218 332 3338 373
rect 3442 373 3478 392
rect 3524 392 3703 419
rect 3524 373 3562 392
rect 3442 332 3562 373
rect 3666 373 3703 392
rect 3749 392 3928 419
rect 3749 373 3786 392
rect 3666 332 3786 373
rect 3890 373 3928 392
rect 3974 392 4147 419
rect 3974 373 4010 392
rect 3890 332 4010 373
rect 4114 373 4147 392
rect 4193 392 4374 419
rect 4193 373 4234 392
rect 4114 332 4234 373
rect 4338 373 4374 392
rect 4420 392 4599 419
rect 4420 373 4458 392
rect 4338 332 4458 373
rect 4562 373 4599 392
rect 4645 392 4824 419
rect 4645 373 4682 392
rect 4562 332 4682 373
rect 4786 373 4824 392
rect 4870 392 5048 419
rect 4870 373 4906 392
rect 4786 332 4906 373
rect 5010 373 5048 392
rect 5094 392 5270 419
rect 5094 373 5130 392
rect 5010 332 5130 373
rect 5234 373 5270 392
rect 5316 392 5498 419
rect 5316 373 5354 392
rect 5234 332 5354 373
rect 5458 373 5498 392
rect 5544 392 6250 419
rect 5544 373 5578 392
rect 5458 332 5578 373
rect 5682 332 5802 392
rect 5906 332 6026 392
rect 6130 332 6250 392
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 978 24 1098 68
rect 1202 24 1322 68
rect 1426 24 1546 68
rect 1650 24 1770 68
rect 1874 24 1994 68
rect 2098 24 2218 68
rect 2322 24 2442 68
rect 2546 24 2666 68
rect 2770 24 2890 68
rect 2994 24 3114 68
rect 3218 24 3338 68
rect 3442 24 3562 68
rect 3666 24 3786 68
rect 3890 24 4010 68
rect 4114 24 4234 68
rect 4338 24 4458 68
rect 4562 24 4682 68
rect 4786 24 4906 68
rect 5010 24 5130 68
rect 5234 24 5354 68
rect 5458 24 5578 68
rect 5682 24 5802 68
rect 5906 24 6026 68
rect 6130 24 6250 68
<< polycontact >>
rect 185 477 231 523
rect 673 494 719 540
rect 361 366 407 412
rect 1085 463 1131 509
rect 1287 463 1333 509
rect 1492 463 1538 509
rect 1695 463 1741 509
rect 1901 463 1947 509
rect 2165 463 2211 509
rect 2369 463 2415 509
rect 2816 494 2862 540
rect 3019 494 3065 540
rect 3223 494 3269 540
rect 3427 494 3473 540
rect 3629 494 3675 540
rect 3833 494 3879 540
rect 4038 494 4084 540
rect 4241 494 4287 540
rect 4447 494 4493 540
rect 4651 494 4697 540
rect 4854 494 4900 540
rect 5058 494 5104 540
rect 5260 494 5306 540
rect 5467 494 5513 540
rect 2783 373 2829 419
rect 3032 373 3078 419
rect 3255 373 3301 419
rect 3478 373 3524 419
rect 3703 373 3749 419
rect 3928 373 3974 419
rect 4147 373 4193 419
rect 4374 373 4420 419
rect 4599 373 4645 419
rect 4824 373 4870 419
rect 5048 373 5094 419
rect 5270 373 5316 419
rect 5498 373 5544 419
<< metal1 >>
rect 0 927 6384 1098
rect 0 920 2711 927
rect 0 918 301 920
rect 347 918 983 920
rect 972 874 983 918
rect 1029 918 1391 920
rect 1029 874 1040 918
rect 1380 874 1391 918
rect 1437 918 1799 920
rect 1437 874 1448 918
rect 1788 874 1799 918
rect 1845 918 2267 920
rect 1845 874 1856 918
rect 2256 874 2267 918
rect 2313 918 2711 920
rect 2313 874 2324 918
rect 2700 881 2711 918
rect 2757 918 3119 927
rect 2757 881 2768 918
rect 3108 881 3119 918
rect 3165 918 3527 927
rect 3165 881 3176 918
rect 3516 881 3527 918
rect 3573 918 3935 927
rect 3573 881 3584 918
rect 3924 881 3935 918
rect 3981 918 4343 927
rect 3981 881 3992 918
rect 4332 881 4343 918
rect 4389 918 4751 927
rect 4389 881 4400 918
rect 4740 881 4751 918
rect 4797 918 5159 927
rect 4797 881 4808 918
rect 5148 881 5159 918
rect 5205 918 5567 927
rect 5205 881 5216 918
rect 5556 881 5567 918
rect 5613 918 5975 927
rect 5613 881 5624 918
rect 301 769 347 780
rect 585 817 2540 828
rect 585 771 1187 817
rect 97 739 143 750
rect 631 725 1187 771
rect 585 689 1187 725
rect 881 677 1187 689
rect 1233 677 1595 817
rect 1641 677 2003 817
rect 2049 770 2540 817
rect 2049 724 2471 770
rect 2517 724 2540 770
rect 2049 677 2540 724
rect 881 666 2540 677
rect 2904 824 5818 835
rect 2904 778 3323 824
rect 2904 732 2915 778
rect 2961 732 3323 778
rect 2904 684 3323 732
rect 3369 684 3731 824
rect 3777 684 4139 824
rect 4185 684 4547 824
rect 4593 684 4955 824
rect 5001 684 5363 824
rect 5409 684 5771 824
rect 5817 684 5818 824
rect 6021 918 6384 927
rect 5975 776 6021 787
rect 2904 673 5818 684
rect 143 599 719 634
rect 97 588 719 599
rect 109 523 315 542
rect 109 477 185 523
rect 231 477 315 523
rect 109 466 315 477
rect 361 412 407 588
rect 673 540 719 588
rect 673 483 719 494
rect 789 632 835 643
rect 789 437 835 586
rect 361 320 407 366
rect 38 274 49 320
rect 95 274 407 320
rect 629 391 835 437
rect 629 298 675 391
rect 881 331 927 666
rect 2471 551 2540 666
rect 1060 509 2425 542
rect 1060 463 1085 509
rect 1131 463 1287 509
rect 1333 463 1492 509
rect 1538 463 1695 509
rect 1741 463 1901 509
rect 1947 463 2165 509
rect 2211 463 2369 509
rect 2415 463 2425 509
rect 2471 540 5524 551
rect 2471 494 2816 540
rect 2862 494 3019 540
rect 3065 494 3223 540
rect 3269 494 3427 540
rect 3473 494 3629 540
rect 3675 494 3833 540
rect 3879 494 4038 540
rect 4084 494 4241 540
rect 4287 494 4447 540
rect 4493 494 4651 540
rect 4697 494 4854 540
rect 4900 494 5058 540
rect 5104 494 5260 540
rect 5306 494 5467 540
rect 5513 494 5524 540
rect 1060 430 2425 463
rect 497 287 675 298
rect 543 217 675 287
rect 721 320 927 331
rect 2771 419 5555 432
rect 2771 373 2783 419
rect 2829 373 3032 419
rect 3078 373 3255 419
rect 3301 373 3478 419
rect 3524 373 3703 419
rect 3749 373 3928 419
rect 3974 373 4147 419
rect 4193 373 4374 419
rect 4420 373 4599 419
rect 4645 373 4824 419
rect 4870 373 5048 419
rect 5094 373 5270 419
rect 5316 373 5498 419
rect 5544 373 5555 419
rect 2771 330 2829 373
rect 767 274 927 320
rect 721 263 927 274
rect 1127 319 2829 330
rect 5706 330 5818 673
rect 5706 327 6101 330
rect 1127 272 1575 319
rect 1173 226 1575 272
rect 1127 217 1575 226
rect 543 179 1575 217
rect 1621 179 2023 319
rect 2069 179 2471 319
rect 2517 179 2829 319
rect 543 173 2829 179
rect 2919 319 6101 327
rect 2919 272 3367 319
rect 2965 226 3367 272
rect 2919 179 3367 226
rect 3413 179 3815 319
rect 3861 179 4263 319
rect 4309 179 4711 319
rect 4757 179 5159 319
rect 5205 179 5607 319
rect 5653 272 6101 319
rect 5653 226 6055 272
rect 5653 179 6101 226
rect 2919 173 6101 179
rect 6279 221 6325 232
rect 543 171 1173 173
rect 273 128 319 139
rect 497 136 543 147
rect 0 82 273 90
rect 854 90 865 125
rect 319 82 865 90
rect 0 79 865 82
rect 911 90 922 125
rect 1340 90 1351 127
rect 911 81 1351 90
rect 1397 90 1408 127
rect 1788 90 1799 127
rect 1397 81 1799 90
rect 1845 90 1856 127
rect 2236 90 2247 127
rect 1845 81 2247 90
rect 2293 90 2304 127
rect 2681 90 2695 127
rect 2293 81 2695 90
rect 2741 90 2756 127
rect 3132 90 3143 127
rect 2741 81 3143 90
rect 3189 90 3200 127
rect 3580 90 3591 127
rect 3189 81 3591 90
rect 3637 90 3648 127
rect 4028 90 4039 127
rect 3637 81 4039 90
rect 4085 90 4096 127
rect 4476 90 4487 127
rect 4085 81 4487 90
rect 4533 90 4544 127
rect 4924 90 4935 127
rect 4533 81 4935 90
rect 4981 90 4992 127
rect 5372 90 5383 127
rect 4981 81 5383 90
rect 5429 90 5440 127
rect 5820 90 5831 127
rect 5429 81 5831 90
rect 5877 90 5888 127
rect 5877 81 6279 90
rect 6325 81 6384 90
rect 911 79 6384 81
rect 0 -90 6384 79
<< labels >>
flabel metal1 s 109 466 315 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1060 430 2425 542 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 6384 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 6279 139 6325 232 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2904 673 5818 835 0 FreeSans 200 0 0 0 Z
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 5706 330 5818 673 1 Z
port 3 nsew default output
rlabel metal1 s 5706 327 6101 330 1 Z
port 3 nsew default output
rlabel metal1 s 2919 173 6101 327 1 Z
port 3 nsew default output
rlabel metal1 s 5975 881 6021 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5556 881 5624 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5148 881 5216 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4740 881 4808 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4332 881 4400 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3924 881 3992 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3516 881 3584 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3108 881 3176 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2700 881 2768 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2256 881 2324 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1788 881 1856 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1380 881 1448 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 972 881 1040 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 881 347 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5975 874 6021 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2256 874 2324 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1788 874 1856 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1380 874 1448 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 972 874 1040 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 874 347 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5975 776 6021 874 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 776 347 874 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 769 347 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6279 127 6325 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6279 125 6325 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5820 125 5888 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5372 125 5440 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4924 125 4992 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4476 125 4544 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4028 125 4096 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3580 125 3648 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 125 3200 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2681 125 2756 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 125 2304 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1788 125 1856 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1340 125 1408 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6279 90 6325 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5820 90 5888 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5372 90 5440 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4924 90 4992 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4476 90 4544 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4028 90 4096 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3580 90 3648 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 90 3200 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2681 90 2756 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 90 2304 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1788 90 1856 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1340 90 1408 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 854 90 922 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 6384 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6384 1008
string GDS_END 1380550
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1367714
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
