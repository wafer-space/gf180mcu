magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< metal1 >>
rect 28753 4280 29077 4292
rect 28753 4228 28765 4280
rect 28817 4228 28889 4280
rect 28941 4228 29013 4280
rect 29065 4228 29077 4280
rect 28753 4156 29077 4228
rect 28753 4104 28765 4156
rect 28817 4104 28889 4156
rect 28941 4104 29013 4156
rect 29065 4104 29077 4156
rect 28753 4032 29077 4104
rect 28753 3980 28765 4032
rect 28817 3980 28889 4032
rect 28941 3980 29013 4032
rect 29065 3980 29077 4032
rect 28753 3908 29077 3980
rect 28753 3856 28765 3908
rect 28817 3856 28889 3908
rect 28941 3856 29013 3908
rect 29065 3856 29077 3908
rect 28753 3844 29077 3856
rect 59890 4280 60214 4292
rect 59890 4228 59902 4280
rect 59954 4228 60026 4280
rect 60078 4228 60150 4280
rect 60202 4228 60214 4280
rect 59890 4156 60214 4228
rect 59890 4104 59902 4156
rect 59954 4104 60026 4156
rect 60078 4104 60150 4156
rect 60202 4104 60214 4156
rect 59890 4032 60214 4104
rect 59890 3980 59902 4032
rect 59954 3980 60026 4032
rect 60078 3980 60150 4032
rect 60202 3980 60214 4032
rect 59890 3908 60214 3980
rect 59890 3856 59902 3908
rect 59954 3856 60026 3908
rect 60078 3856 60150 3908
rect 60202 3856 60214 3908
rect 59890 3844 60214 3856
<< via1 >>
rect 28765 4228 28817 4280
rect 28889 4228 28941 4280
rect 29013 4228 29065 4280
rect 28765 4104 28817 4156
rect 28889 4104 28941 4156
rect 29013 4104 29065 4156
rect 28765 3980 28817 4032
rect 28889 3980 28941 4032
rect 29013 3980 29065 4032
rect 28765 3856 28817 3908
rect 28889 3856 28941 3908
rect 29013 3856 29065 3908
rect 59902 4228 59954 4280
rect 60026 4228 60078 4280
rect 60150 4228 60202 4280
rect 59902 4104 59954 4156
rect 60026 4104 60078 4156
rect 60150 4104 60202 4156
rect 59902 3980 59954 4032
rect 60026 3980 60078 4032
rect 60150 3980 60202 4032
rect 59902 3856 59954 3908
rect 60026 3856 60078 3908
rect 60150 3856 60202 3908
<< metal2 >>
rect 28753 4282 29077 4292
rect 28753 4226 28763 4282
rect 28819 4226 28887 4282
rect 28943 4226 29011 4282
rect 29067 4226 29077 4282
rect 28753 4158 29077 4226
rect 28753 4102 28763 4158
rect 28819 4102 28887 4158
rect 28943 4102 29011 4158
rect 29067 4102 29077 4158
rect 28753 4034 29077 4102
rect 28753 3978 28763 4034
rect 28819 3978 28887 4034
rect 28943 3978 29011 4034
rect 29067 3978 29077 4034
rect 28753 3910 29077 3978
rect 28753 3854 28763 3910
rect 28819 3854 28887 3910
rect 28943 3854 29011 3910
rect 29067 3854 29077 3910
rect 28753 3844 29077 3854
rect 59830 4282 60272 6104
rect 59830 4226 59900 4282
rect 59956 4226 60024 4282
rect 60080 4226 60148 4282
rect 60204 4226 60272 4282
rect 59830 4158 60272 4226
rect 59830 4102 59900 4158
rect 59956 4102 60024 4158
rect 60080 4102 60148 4158
rect 60204 4102 60272 4158
rect 59830 4034 60272 4102
rect 59830 3978 59900 4034
rect 59956 3978 60024 4034
rect 60080 3978 60148 4034
rect 60204 3978 60272 4034
rect 59830 3910 60272 3978
rect 59830 3854 59900 3910
rect 59956 3854 60024 3910
rect 60080 3854 60148 3910
rect 60204 3854 60272 3910
rect 59830 3357 60272 3854
<< via2 >>
rect 28763 4280 28819 4282
rect 28763 4228 28765 4280
rect 28765 4228 28817 4280
rect 28817 4228 28819 4280
rect 28763 4226 28819 4228
rect 28887 4280 28943 4282
rect 28887 4228 28889 4280
rect 28889 4228 28941 4280
rect 28941 4228 28943 4280
rect 28887 4226 28943 4228
rect 29011 4280 29067 4282
rect 29011 4228 29013 4280
rect 29013 4228 29065 4280
rect 29065 4228 29067 4280
rect 29011 4226 29067 4228
rect 28763 4156 28819 4158
rect 28763 4104 28765 4156
rect 28765 4104 28817 4156
rect 28817 4104 28819 4156
rect 28763 4102 28819 4104
rect 28887 4156 28943 4158
rect 28887 4104 28889 4156
rect 28889 4104 28941 4156
rect 28941 4104 28943 4156
rect 28887 4102 28943 4104
rect 29011 4156 29067 4158
rect 29011 4104 29013 4156
rect 29013 4104 29065 4156
rect 29065 4104 29067 4156
rect 29011 4102 29067 4104
rect 28763 4032 28819 4034
rect 28763 3980 28765 4032
rect 28765 3980 28817 4032
rect 28817 3980 28819 4032
rect 28763 3978 28819 3980
rect 28887 4032 28943 4034
rect 28887 3980 28889 4032
rect 28889 3980 28941 4032
rect 28941 3980 28943 4032
rect 28887 3978 28943 3980
rect 29011 4032 29067 4034
rect 29011 3980 29013 4032
rect 29013 3980 29065 4032
rect 29065 3980 29067 4032
rect 29011 3978 29067 3980
rect 28763 3908 28819 3910
rect 28763 3856 28765 3908
rect 28765 3856 28817 3908
rect 28817 3856 28819 3908
rect 28763 3854 28819 3856
rect 28887 3908 28943 3910
rect 28887 3856 28889 3908
rect 28889 3856 28941 3908
rect 28941 3856 28943 3908
rect 28887 3854 28943 3856
rect 29011 3908 29067 3910
rect 29011 3856 29013 3908
rect 29013 3856 29065 3908
rect 29065 3856 29067 3908
rect 29011 3854 29067 3856
rect 59900 4280 59956 4282
rect 59900 4228 59902 4280
rect 59902 4228 59954 4280
rect 59954 4228 59956 4280
rect 59900 4226 59956 4228
rect 60024 4280 60080 4282
rect 60024 4228 60026 4280
rect 60026 4228 60078 4280
rect 60078 4228 60080 4280
rect 60024 4226 60080 4228
rect 60148 4280 60204 4282
rect 60148 4228 60150 4280
rect 60150 4228 60202 4280
rect 60202 4228 60204 4280
rect 60148 4226 60204 4228
rect 59900 4156 59956 4158
rect 59900 4104 59902 4156
rect 59902 4104 59954 4156
rect 59954 4104 59956 4156
rect 59900 4102 59956 4104
rect 60024 4156 60080 4158
rect 60024 4104 60026 4156
rect 60026 4104 60078 4156
rect 60078 4104 60080 4156
rect 60024 4102 60080 4104
rect 60148 4156 60204 4158
rect 60148 4104 60150 4156
rect 60150 4104 60202 4156
rect 60202 4104 60204 4156
rect 60148 4102 60204 4104
rect 59900 4032 59956 4034
rect 59900 3980 59902 4032
rect 59902 3980 59954 4032
rect 59954 3980 59956 4032
rect 59900 3978 59956 3980
rect 60024 4032 60080 4034
rect 60024 3980 60026 4032
rect 60026 3980 60078 4032
rect 60078 3980 60080 4032
rect 60024 3978 60080 3980
rect 60148 4032 60204 4034
rect 60148 3980 60150 4032
rect 60150 3980 60202 4032
rect 60202 3980 60204 4032
rect 60148 3978 60204 3980
rect 59900 3908 59956 3910
rect 59900 3856 59902 3908
rect 59902 3856 59954 3908
rect 59954 3856 59956 3908
rect 59900 3854 59956 3856
rect 60024 3908 60080 3910
rect 60024 3856 60026 3908
rect 60026 3856 60078 3908
rect 60078 3856 60080 3908
rect 60024 3854 60080 3856
rect 60148 3908 60204 3910
rect 60148 3856 60150 3908
rect 60150 3856 60202 3908
rect 60202 3856 60204 3908
rect 60148 3854 60204 3856
<< metal3 >>
rect 28753 4282 29077 4292
rect 28753 4226 28763 4282
rect 28819 4226 28887 4282
rect 28943 4226 29011 4282
rect 29067 4226 29077 4282
rect 28753 4158 29077 4226
rect 28753 4102 28763 4158
rect 28819 4102 28887 4158
rect 28943 4102 29011 4158
rect 29067 4102 29077 4158
rect 28753 4034 29077 4102
rect 28753 3978 28763 4034
rect 28819 3978 28887 4034
rect 28943 3978 29011 4034
rect 29067 3978 29077 4034
rect 28753 3910 29077 3978
rect 28753 3854 28763 3910
rect 28819 3854 28887 3910
rect 28943 3854 29011 3910
rect 29067 3854 29077 3910
rect 28753 3844 29077 3854
rect 59890 4282 60214 4292
rect 59890 4226 59900 4282
rect 59956 4226 60024 4282
rect 60080 4226 60148 4282
rect 60204 4226 60214 4282
rect 59890 4158 60214 4226
rect 59890 4102 59900 4158
rect 59956 4102 60024 4158
rect 60080 4102 60148 4158
rect 60204 4102 60214 4158
rect 59890 4034 60214 4102
rect 59890 3978 59900 4034
rect 59956 3978 60024 4034
rect 60080 3978 60148 4034
rect 60204 3978 60214 4034
rect 59890 3910 60214 3978
rect 59890 3854 59900 3910
rect 59956 3854 60024 3910
rect 60080 3854 60148 3910
rect 60204 3854 60214 3910
rect 59890 3844 60214 3854
use M2_M14310590878169_256x8m81  M2_M14310590878169_256x8m81_0
timestamp 1755724134
transform 1 0 60052 0 1 4068
box 0 0 1 1
use M2_M14310590878169_256x8m81  M2_M14310590878169_256x8m81_1
timestamp 1755724134
transform 1 0 28915 0 1 4068
box 0 0 1 1
use M3_M24310590878170_256x8m81  M3_M24310590878170_256x8m81_0
timestamp 1755724134
transform 1 0 60052 0 1 4068
box 0 0 1 1
use M3_M24310590878170_256x8m81  M3_M24310590878170_256x8m81_1
timestamp 1755724134
transform 1 0 28915 0 1 4068
box 0 0 1 1
use power_route_01_256x8m81  power_route_01_256x8m81_0
timestamp 1755724134
transform -1 0 25893 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_1
timestamp 1755724134
transform 1 0 9233 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_2
timestamp 1755724134
transform 1 0 20033 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_3
timestamp 1755724134
transform 1 0 14633 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_4
timestamp 1755724134
transform 1 0 63409 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_5
timestamp 1755724134
transform 1 0 79609 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_6
timestamp 1755724134
transform 1 0 74209 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_7
timestamp 1755724134
transform 1 0 68810 0 1 67814
box -511 0 1714 2425
use power_route_01_256x8m81  power_route_01_256x8m81_8
timestamp 1755724134
transform 1 0 3833 0 1 67814
box -511 0 1714 2425
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_0
timestamp 1755724134
transform 1 0 -1418 0 1 65089
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_1
timestamp 1755724134
transform 1 0 -1418 0 1 61489
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_2
timestamp 1755724134
transform 1 0 -1418 0 1 63289
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_3
timestamp 1755724134
transform 1 0 -1418 0 1 54289
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_4
timestamp 1755724134
transform 1 0 -1418 0 1 56089
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_5
timestamp 1755724134
transform 1 0 -1418 0 1 59689
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_6
timestamp 1755724134
transform 1 0 -1418 0 1 57889
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_7
timestamp 1755724134
transform 1 0 -1418 0 1 52489
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_8
timestamp 1755724134
transform 1 0 -1418 0 1 50689
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_9
timestamp 1755724134
transform 1 0 -1418 0 1 47089
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_10
timestamp 1755724134
transform 1 0 -1418 0 1 48889
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_11
timestamp 1755724134
transform 1 0 -1418 0 1 39889
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_12
timestamp 1755724134
transform 1 0 -1418 0 1 41689
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_13
timestamp 1755724134
transform 1 0 -1418 0 1 45289
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_14
timestamp 1755724134
transform 1 0 -1418 0 1 43489
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_15
timestamp 1755724134
transform 1 0 -1418 0 1 38089
box 3339 -250 30611 1350
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_16
timestamp 1755724134
transform 1 0 -1418 0 1 66889
box 3339 -250 30611 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_0
timestamp 1755724134
transform -1 0 91632 0 1 39889
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_1
timestamp 1755724134
transform -1 0 91632 0 1 41689
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_2
timestamp 1755724134
transform -1 0 91632 0 1 43489
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_3
timestamp 1755724134
transform -1 0 91632 0 1 45289
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_4
timestamp 1755724134
transform -1 0 91632 0 1 47089
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_5
timestamp 1755724134
transform -1 0 91632 0 1 48889
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_6
timestamp 1755724134
transform -1 0 91632 0 1 50689
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_7
timestamp 1755724134
transform -1 0 91632 0 1 52489
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_8
timestamp 1755724134
transform -1 0 91632 0 1 54289
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_9
timestamp 1755724134
transform -1 0 91632 0 1 56089
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_10
timestamp 1755724134
transform -1 0 91632 0 1 57889
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_11
timestamp 1755724134
transform -1 0 91632 0 1 59689
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_12
timestamp 1755724134
transform -1 0 91632 0 1 61489
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_13
timestamp 1755724134
transform -1 0 91632 0 1 63289
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_14
timestamp 1755724134
transform -1 0 91632 0 1 65089
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_15
timestamp 1755724134
transform -1 0 91632 0 1 66889
box 3339 -250 29240 1350
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_16
timestamp 1755724134
transform -1 0 91632 0 1 38089
box 3339 -250 29240 1350
use power_route_04_256x8m81  power_route_04_256x8m81_0
timestamp 1755724134
transform -1 0 91632 0 1 244
box 3339 2101 6632 52645
use power_route_04_256x8m81  power_route_04_256x8m81_1
timestamp 1755724134
transform 1 0 -1418 0 1 244
box 3339 2101 6632 52645
use power_route_05_256x8m81  power_route_05_256x8m81_0
timestamp 1755724134
transform 1 0 19656 0 1 230
box -8 2115 1235 7462
use power_route_05_256x8m81  power_route_05_256x8m81_1
timestamp 1755724134
transform 1 0 68431 0 1 230
box -8 2115 1235 7462
use power_route_05_256x8m81  power_route_05_256x8m81_2
timestamp 1755724134
transform 1 0 79230 0 1 230
box -8 2115 1235 7462
use power_route_05_256x8m81  power_route_05_256x8m81_3
timestamp 1755724134
transform 1 0 8856 0 1 230
box -8 2115 1235 7462
use power_route_06_256x8m81  power_route_06_256x8m81_0
timestamp 1755724134
transform 1 0 61241 0 1 230
box -7 2115 1234 18431
use power_route_06_256x8m81  power_route_06_256x8m81_1
timestamp 1755724134
transform 1 0 26784 0 1 230
box -7 2115 1234 18431
use power_route_07_256x8m81  power_route_07_256x8m81_0
timestamp 1755724134
transform 1 0 40746 0 1 230
box -8 3065 1235 7462
use power_route_07_256x8m81  power_route_07_256x8m81_1
timestamp 1755724134
transform 1 0 38926 0 1 230
box -8 3065 1235 7462
<< properties >>
string GDS_END 2395660
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2392430
<< end >>
