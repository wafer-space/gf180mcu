magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1755724134
transform 1 0 4563 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1755724134
transform 1 0 3891 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1755724134
transform 1 0 400 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1755724134
transform 1 0 1520 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1755724134
transform 1 0 5749 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1755724134
transform 1 0 5973 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1755724134
transform 1 0 1072 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_7
timestamp 1755724134
transform 1 0 848 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_8
timestamp 1755724134
transform 1 0 4787 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_9
timestamp 1755724134
transform 1 0 3667 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_10
timestamp 1755724134
transform 1 0 5525 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_11
timestamp 1755724134
transform 1 0 6197 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_12
timestamp 1755724134
transform 1 0 2929 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_13
timestamp 1755724134
transform 1 0 2257 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_14
timestamp 1755724134
transform 1 0 2705 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_15
timestamp 1755724134
transform 1 0 2481 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_16
timestamp 1755724134
transform 1 0 6421 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_17
timestamp 1755724134
transform 1 0 3153 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_18
timestamp 1755724134
transform 1 0 2033 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_19
timestamp 1755724134
transform 1 0 5301 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_20
timestamp 1755724134
transform 1 0 1296 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_21
timestamp 1755724134
transform 1 0 624 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_22
timestamp 1755724134
transform 1 0 4115 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_23
timestamp 1755724134
transform 1 0 4339 0 1 2018
box 0 0 1 1
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_0
timestamp 1755724134
transform 1 0 2594 0 1 1002
box 0 0 1 1
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_1
timestamp 1755724134
transform 1 0 4227 0 1 1002
box 0 0 1 1
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_2
timestamp 1755724134
transform 1 0 5861 0 1 1002
box 0 0 1 1
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_3
timestamp 1755724134
transform 1 0 960 0 1 1002
box 0 0 1 1
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_0
timestamp 1755724134
transform 1 0 960 0 1 1002
box 0 0 1 1
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_1
timestamp 1755724134
transform 1 0 4227 0 1 1002
box 0 0 1 1
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_2
timestamp 1755724134
transform 1 0 5861 0 1 1002
box 0 0 1 1
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_3
timestamp 1755724134
transform 1 0 2594 0 1 1002
box 0 0 1 1
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_0
timestamp 1755724134
transform -1 0 4372 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_1
timestamp 1755724134
transform -1 0 6006 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_2
timestamp 1755724134
transform -1 0 2738 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_3
timestamp 1755724134
transform -1 0 1105 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_4
timestamp 1755724134
transform 1 0 4082 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_5
timestamp 1755724134
transform 1 0 5716 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_6
timestamp 1755724134
transform 1 0 2448 0 1 7069
box 145 -5906 818 -136
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_7
timestamp 1755724134
transform 1 0 815 0 1 7069
box 145 -5906 818 -136
<< properties >>
string GDS_END 967942
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 965850
<< end >>
