magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 758 870
<< pwell >>
rect -86 -86 758 352
<< metal1 >>
rect 0 724 672 844
rect 262 603 330 724
rect 141 348 318 430
rect 141 207 216 348
rect 513 321 586 664
rect 262 60 330 185
rect 468 113 586 321
rect 0 -60 672 60
<< obsm1 >>
rect 49 551 115 676
rect 49 504 454 551
rect 49 113 95 504
rect 386 376 454 504
<< labels >>
rlabel metal1 s 141 207 216 348 6 I
port 1 nsew default input
rlabel metal1 s 141 348 318 430 6 I
port 1 nsew default input
rlabel metal1 s 468 113 586 321 6 Z
port 2 nsew default output
rlabel metal1 s 513 321 586 664 6 Z
port 2 nsew default output
rlabel metal1 s 262 603 330 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 672 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 758 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 758 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 672 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 185 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1443700
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1441056
<< end >>
