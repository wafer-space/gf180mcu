magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< metal1 >>
rect 1398 956 1578 968
rect 1398 904 1410 956
rect 1566 904 1578 956
rect 1398 892 1578 904
rect 1818 959 2608 971
rect 1818 803 1830 959
rect 1882 809 2608 959
rect 2784 968 2860 980
rect 2784 812 2796 968
rect 2848 812 2860 968
rect 1882 803 1894 809
rect 1818 791 1894 803
rect 2784 800 2860 812
rect 2900 -489 2976 -477
rect 2900 -645 2912 -489
rect 2964 -645 2976 -489
rect 1299 -1157 1375 -1145
rect 1299 -1313 1311 -1157
rect 1363 -1313 1375 -1157
rect 1299 -1325 1375 -1313
rect 2900 -2007 2976 -645
rect 2282 -2083 2976 -2007
<< via1 >>
rect 1410 904 1566 956
rect 1830 803 1882 959
rect 2796 812 2848 968
rect 2912 -645 2964 -489
rect 1311 -1313 1363 -1157
<< metal2 >>
rect 1206 1153 1894 1229
rect 1206 -967 1282 1153
rect 1502 968 1578 980
rect 1398 956 1578 968
rect 1398 904 1410 956
rect 1566 904 1578 956
rect 1398 892 1578 904
rect 1148 -1043 1282 -967
rect 1148 -1426 1224 -1043
rect 1502 -1145 1578 892
rect 1818 959 1894 1153
rect 1818 803 1830 959
rect 1882 803 1894 959
rect 1818 791 1894 803
rect 2784 968 2860 981
rect 2784 812 2796 968
rect 2848 812 2860 968
rect 2784 -477 2860 812
rect 2784 -489 2976 -477
rect 2784 -553 2912 -489
rect 2900 -645 2912 -553
rect 2964 -645 2976 -489
rect 2900 -657 2976 -645
rect 1299 -1157 1578 -1145
rect 1299 -1313 1311 -1157
rect 1363 -1221 1578 -1157
rect 1363 -1313 1375 -1221
rect 1299 -1325 1375 -1313
rect 1148 -1493 1339 -1426
rect 1263 -1611 1339 -1493
use comp018green_std_nand2  comp018green_std_nand2_0
timestamp 1755724134
transform 1 0 2168 0 -1 2153
box -83 11 1139 2586
use comp018green_std_nand2  comp018green_std_nand2_1
timestamp 1755724134
transform 1 0 1202 0 -1 2153
box -83 11 1139 2586
use comp018green_std_xor2  comp018green_std_xor2_0
timestamp 1755724134
transform 1 0 511 0 1 -3277
box -83 0 2361 2575
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1755724134
transform 0 1 1488 1 0 930
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1755724134
transform 1 0 1856 0 -1 881
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1755724134
transform 1 0 2822 0 -1 890
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1755724134
transform 1 0 2938 0 1 -567
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1755724134
transform 1 0 1337 0 1 -1235
box 0 0 1 1
<< labels >>
rlabel metal2 s 2185 -2041 2185 -2041 4 PD_IN
port 1 nsew
rlabel metal1 s 1861 1095 1861 1095 4 PUB_OUT
port 2 nsew
rlabel metal1 s 2840 1095 2840 1095 4 PDB_OUT
port 3 nsew
rlabel metal1 s 781 -825 781 -825 4 VDD
port 4 nsew
rlabel metal1 s 755 -3232 755 -3232 4 VSS
port 5 nsew
<< properties >>
string GDS_END 1532816
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1531596
string path 57.050 -51.125 73.450 -51.125 73.450 -11.925 
<< end >>
