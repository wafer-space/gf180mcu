magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< deepnwell >>
rect -680 -680 2680 2680
<< pbase >>
rect -180 -180 2180 2180
<< ndiff >>
rect 0 1923 2000 2000
rect 0 1877 77 1923
rect 123 1877 197 1923
rect 243 1877 317 1923
rect 363 1877 437 1923
rect 483 1877 557 1923
rect 603 1877 677 1923
rect 723 1877 797 1923
rect 843 1877 917 1923
rect 963 1877 1037 1923
rect 1083 1877 1157 1923
rect 1203 1877 1277 1923
rect 1323 1877 1397 1923
rect 1443 1877 1517 1923
rect 1563 1877 1637 1923
rect 1683 1877 1757 1923
rect 1803 1877 1877 1923
rect 1923 1877 2000 1923
rect 0 1803 2000 1877
rect 0 1757 77 1803
rect 123 1757 197 1803
rect 243 1757 317 1803
rect 363 1757 437 1803
rect 483 1757 557 1803
rect 603 1757 677 1803
rect 723 1757 797 1803
rect 843 1757 917 1803
rect 963 1757 1037 1803
rect 1083 1757 1157 1803
rect 1203 1757 1277 1803
rect 1323 1757 1397 1803
rect 1443 1757 1517 1803
rect 1563 1757 1637 1803
rect 1683 1757 1757 1803
rect 1803 1757 1877 1803
rect 1923 1757 2000 1803
rect 0 1683 2000 1757
rect 0 1637 77 1683
rect 123 1637 197 1683
rect 243 1637 317 1683
rect 363 1637 437 1683
rect 483 1637 557 1683
rect 603 1637 677 1683
rect 723 1637 797 1683
rect 843 1637 917 1683
rect 963 1637 1037 1683
rect 1083 1637 1157 1683
rect 1203 1637 1277 1683
rect 1323 1637 1397 1683
rect 1443 1637 1517 1683
rect 1563 1637 1637 1683
rect 1683 1637 1757 1683
rect 1803 1637 1877 1683
rect 1923 1637 2000 1683
rect 0 1563 2000 1637
rect 0 1517 77 1563
rect 123 1517 197 1563
rect 243 1517 317 1563
rect 363 1517 437 1563
rect 483 1517 557 1563
rect 603 1517 677 1563
rect 723 1517 797 1563
rect 843 1517 917 1563
rect 963 1517 1037 1563
rect 1083 1517 1157 1563
rect 1203 1517 1277 1563
rect 1323 1517 1397 1563
rect 1443 1517 1517 1563
rect 1563 1517 1637 1563
rect 1683 1517 1757 1563
rect 1803 1517 1877 1563
rect 1923 1517 2000 1563
rect 0 1443 2000 1517
rect 0 1397 77 1443
rect 123 1397 197 1443
rect 243 1397 317 1443
rect 363 1397 437 1443
rect 483 1397 557 1443
rect 603 1397 677 1443
rect 723 1397 797 1443
rect 843 1397 917 1443
rect 963 1397 1037 1443
rect 1083 1397 1157 1443
rect 1203 1397 1277 1443
rect 1323 1397 1397 1443
rect 1443 1397 1517 1443
rect 1563 1397 1637 1443
rect 1683 1397 1757 1443
rect 1803 1397 1877 1443
rect 1923 1397 2000 1443
rect 0 1323 2000 1397
rect 0 1277 77 1323
rect 123 1277 197 1323
rect 243 1277 317 1323
rect 363 1277 437 1323
rect 483 1277 557 1323
rect 603 1277 677 1323
rect 723 1277 797 1323
rect 843 1277 917 1323
rect 963 1277 1037 1323
rect 1083 1277 1157 1323
rect 1203 1277 1277 1323
rect 1323 1277 1397 1323
rect 1443 1277 1517 1323
rect 1563 1277 1637 1323
rect 1683 1277 1757 1323
rect 1803 1277 1877 1323
rect 1923 1277 2000 1323
rect 0 1203 2000 1277
rect 0 1157 77 1203
rect 123 1157 197 1203
rect 243 1157 317 1203
rect 363 1157 437 1203
rect 483 1157 557 1203
rect 603 1157 677 1203
rect 723 1157 797 1203
rect 843 1157 917 1203
rect 963 1157 1037 1203
rect 1083 1157 1157 1203
rect 1203 1157 1277 1203
rect 1323 1157 1397 1203
rect 1443 1157 1517 1203
rect 1563 1157 1637 1203
rect 1683 1157 1757 1203
rect 1803 1157 1877 1203
rect 1923 1157 2000 1203
rect 0 1083 2000 1157
rect 0 1037 77 1083
rect 123 1037 197 1083
rect 243 1037 317 1083
rect 363 1037 437 1083
rect 483 1037 557 1083
rect 603 1037 677 1083
rect 723 1037 797 1083
rect 843 1037 917 1083
rect 963 1037 1037 1083
rect 1083 1037 1157 1083
rect 1203 1037 1277 1083
rect 1323 1037 1397 1083
rect 1443 1037 1517 1083
rect 1563 1037 1637 1083
rect 1683 1037 1757 1083
rect 1803 1037 1877 1083
rect 1923 1037 2000 1083
rect 0 963 2000 1037
rect 0 917 77 963
rect 123 917 197 963
rect 243 917 317 963
rect 363 917 437 963
rect 483 917 557 963
rect 603 917 677 963
rect 723 917 797 963
rect 843 917 917 963
rect 963 917 1037 963
rect 1083 917 1157 963
rect 1203 917 1277 963
rect 1323 917 1397 963
rect 1443 917 1517 963
rect 1563 917 1637 963
rect 1683 917 1757 963
rect 1803 917 1877 963
rect 1923 917 2000 963
rect 0 843 2000 917
rect 0 797 77 843
rect 123 797 197 843
rect 243 797 317 843
rect 363 797 437 843
rect 483 797 557 843
rect 603 797 677 843
rect 723 797 797 843
rect 843 797 917 843
rect 963 797 1037 843
rect 1083 797 1157 843
rect 1203 797 1277 843
rect 1323 797 1397 843
rect 1443 797 1517 843
rect 1563 797 1637 843
rect 1683 797 1757 843
rect 1803 797 1877 843
rect 1923 797 2000 843
rect 0 723 2000 797
rect 0 677 77 723
rect 123 677 197 723
rect 243 677 317 723
rect 363 677 437 723
rect 483 677 557 723
rect 603 677 677 723
rect 723 677 797 723
rect 843 677 917 723
rect 963 677 1037 723
rect 1083 677 1157 723
rect 1203 677 1277 723
rect 1323 677 1397 723
rect 1443 677 1517 723
rect 1563 677 1637 723
rect 1683 677 1757 723
rect 1803 677 1877 723
rect 1923 677 2000 723
rect 0 603 2000 677
rect 0 557 77 603
rect 123 557 197 603
rect 243 557 317 603
rect 363 557 437 603
rect 483 557 557 603
rect 603 557 677 603
rect 723 557 797 603
rect 843 557 917 603
rect 963 557 1037 603
rect 1083 557 1157 603
rect 1203 557 1277 603
rect 1323 557 1397 603
rect 1443 557 1517 603
rect 1563 557 1637 603
rect 1683 557 1757 603
rect 1803 557 1877 603
rect 1923 557 2000 603
rect 0 483 2000 557
rect 0 437 77 483
rect 123 437 197 483
rect 243 437 317 483
rect 363 437 437 483
rect 483 437 557 483
rect 603 437 677 483
rect 723 437 797 483
rect 843 437 917 483
rect 963 437 1037 483
rect 1083 437 1157 483
rect 1203 437 1277 483
rect 1323 437 1397 483
rect 1443 437 1517 483
rect 1563 437 1637 483
rect 1683 437 1757 483
rect 1803 437 1877 483
rect 1923 437 2000 483
rect 0 363 2000 437
rect 0 317 77 363
rect 123 317 197 363
rect 243 317 317 363
rect 363 317 437 363
rect 483 317 557 363
rect 603 317 677 363
rect 723 317 797 363
rect 843 317 917 363
rect 963 317 1037 363
rect 1083 317 1157 363
rect 1203 317 1277 363
rect 1323 317 1397 363
rect 1443 317 1517 363
rect 1563 317 1637 363
rect 1683 317 1757 363
rect 1803 317 1877 363
rect 1923 317 2000 363
rect 0 243 2000 317
rect 0 197 77 243
rect 123 197 197 243
rect 243 197 317 243
rect 363 197 437 243
rect 483 197 557 243
rect 603 197 677 243
rect 723 197 797 243
rect 843 197 917 243
rect 963 197 1037 243
rect 1083 197 1157 243
rect 1203 197 1277 243
rect 1323 197 1397 243
rect 1443 197 1517 243
rect 1563 197 1637 243
rect 1683 197 1757 243
rect 1803 197 1877 243
rect 1923 197 2000 243
rect 0 123 2000 197
rect 0 77 77 123
rect 123 77 197 123
rect 243 77 317 123
rect 363 77 437 123
rect 483 77 557 123
rect 603 77 677 123
rect 723 77 797 123
rect 843 77 917 123
rect 963 77 1037 123
rect 1083 77 1157 123
rect 1203 77 1277 123
rect 1323 77 1397 123
rect 1443 77 1517 123
rect 1563 77 1637 123
rect 1683 77 1757 123
rect 1803 77 1877 123
rect 1923 77 2000 123
rect 0 0 2000 77
<< ndiffc >>
rect 77 1877 123 1923
rect 197 1877 243 1923
rect 317 1877 363 1923
rect 437 1877 483 1923
rect 557 1877 603 1923
rect 677 1877 723 1923
rect 797 1877 843 1923
rect 917 1877 963 1923
rect 1037 1877 1083 1923
rect 1157 1877 1203 1923
rect 1277 1877 1323 1923
rect 1397 1877 1443 1923
rect 1517 1877 1563 1923
rect 1637 1877 1683 1923
rect 1757 1877 1803 1923
rect 1877 1877 1923 1923
rect 77 1757 123 1803
rect 197 1757 243 1803
rect 317 1757 363 1803
rect 437 1757 483 1803
rect 557 1757 603 1803
rect 677 1757 723 1803
rect 797 1757 843 1803
rect 917 1757 963 1803
rect 1037 1757 1083 1803
rect 1157 1757 1203 1803
rect 1277 1757 1323 1803
rect 1397 1757 1443 1803
rect 1517 1757 1563 1803
rect 1637 1757 1683 1803
rect 1757 1757 1803 1803
rect 1877 1757 1923 1803
rect 77 1637 123 1683
rect 197 1637 243 1683
rect 317 1637 363 1683
rect 437 1637 483 1683
rect 557 1637 603 1683
rect 677 1637 723 1683
rect 797 1637 843 1683
rect 917 1637 963 1683
rect 1037 1637 1083 1683
rect 1157 1637 1203 1683
rect 1277 1637 1323 1683
rect 1397 1637 1443 1683
rect 1517 1637 1563 1683
rect 1637 1637 1683 1683
rect 1757 1637 1803 1683
rect 1877 1637 1923 1683
rect 77 1517 123 1563
rect 197 1517 243 1563
rect 317 1517 363 1563
rect 437 1517 483 1563
rect 557 1517 603 1563
rect 677 1517 723 1563
rect 797 1517 843 1563
rect 917 1517 963 1563
rect 1037 1517 1083 1563
rect 1157 1517 1203 1563
rect 1277 1517 1323 1563
rect 1397 1517 1443 1563
rect 1517 1517 1563 1563
rect 1637 1517 1683 1563
rect 1757 1517 1803 1563
rect 1877 1517 1923 1563
rect 77 1397 123 1443
rect 197 1397 243 1443
rect 317 1397 363 1443
rect 437 1397 483 1443
rect 557 1397 603 1443
rect 677 1397 723 1443
rect 797 1397 843 1443
rect 917 1397 963 1443
rect 1037 1397 1083 1443
rect 1157 1397 1203 1443
rect 1277 1397 1323 1443
rect 1397 1397 1443 1443
rect 1517 1397 1563 1443
rect 1637 1397 1683 1443
rect 1757 1397 1803 1443
rect 1877 1397 1923 1443
rect 77 1277 123 1323
rect 197 1277 243 1323
rect 317 1277 363 1323
rect 437 1277 483 1323
rect 557 1277 603 1323
rect 677 1277 723 1323
rect 797 1277 843 1323
rect 917 1277 963 1323
rect 1037 1277 1083 1323
rect 1157 1277 1203 1323
rect 1277 1277 1323 1323
rect 1397 1277 1443 1323
rect 1517 1277 1563 1323
rect 1637 1277 1683 1323
rect 1757 1277 1803 1323
rect 1877 1277 1923 1323
rect 77 1157 123 1203
rect 197 1157 243 1203
rect 317 1157 363 1203
rect 437 1157 483 1203
rect 557 1157 603 1203
rect 677 1157 723 1203
rect 797 1157 843 1203
rect 917 1157 963 1203
rect 1037 1157 1083 1203
rect 1157 1157 1203 1203
rect 1277 1157 1323 1203
rect 1397 1157 1443 1203
rect 1517 1157 1563 1203
rect 1637 1157 1683 1203
rect 1757 1157 1803 1203
rect 1877 1157 1923 1203
rect 77 1037 123 1083
rect 197 1037 243 1083
rect 317 1037 363 1083
rect 437 1037 483 1083
rect 557 1037 603 1083
rect 677 1037 723 1083
rect 797 1037 843 1083
rect 917 1037 963 1083
rect 1037 1037 1083 1083
rect 1157 1037 1203 1083
rect 1277 1037 1323 1083
rect 1397 1037 1443 1083
rect 1517 1037 1563 1083
rect 1637 1037 1683 1083
rect 1757 1037 1803 1083
rect 1877 1037 1923 1083
rect 77 917 123 963
rect 197 917 243 963
rect 317 917 363 963
rect 437 917 483 963
rect 557 917 603 963
rect 677 917 723 963
rect 797 917 843 963
rect 917 917 963 963
rect 1037 917 1083 963
rect 1157 917 1203 963
rect 1277 917 1323 963
rect 1397 917 1443 963
rect 1517 917 1563 963
rect 1637 917 1683 963
rect 1757 917 1803 963
rect 1877 917 1923 963
rect 77 797 123 843
rect 197 797 243 843
rect 317 797 363 843
rect 437 797 483 843
rect 557 797 603 843
rect 677 797 723 843
rect 797 797 843 843
rect 917 797 963 843
rect 1037 797 1083 843
rect 1157 797 1203 843
rect 1277 797 1323 843
rect 1397 797 1443 843
rect 1517 797 1563 843
rect 1637 797 1683 843
rect 1757 797 1803 843
rect 1877 797 1923 843
rect 77 677 123 723
rect 197 677 243 723
rect 317 677 363 723
rect 437 677 483 723
rect 557 677 603 723
rect 677 677 723 723
rect 797 677 843 723
rect 917 677 963 723
rect 1037 677 1083 723
rect 1157 677 1203 723
rect 1277 677 1323 723
rect 1397 677 1443 723
rect 1517 677 1563 723
rect 1637 677 1683 723
rect 1757 677 1803 723
rect 1877 677 1923 723
rect 77 557 123 603
rect 197 557 243 603
rect 317 557 363 603
rect 437 557 483 603
rect 557 557 603 603
rect 677 557 723 603
rect 797 557 843 603
rect 917 557 963 603
rect 1037 557 1083 603
rect 1157 557 1203 603
rect 1277 557 1323 603
rect 1397 557 1443 603
rect 1517 557 1563 603
rect 1637 557 1683 603
rect 1757 557 1803 603
rect 1877 557 1923 603
rect 77 437 123 483
rect 197 437 243 483
rect 317 437 363 483
rect 437 437 483 483
rect 557 437 603 483
rect 677 437 723 483
rect 797 437 843 483
rect 917 437 963 483
rect 1037 437 1083 483
rect 1157 437 1203 483
rect 1277 437 1323 483
rect 1397 437 1443 483
rect 1517 437 1563 483
rect 1637 437 1683 483
rect 1757 437 1803 483
rect 1877 437 1923 483
rect 77 317 123 363
rect 197 317 243 363
rect 317 317 363 363
rect 437 317 483 363
rect 557 317 603 363
rect 677 317 723 363
rect 797 317 843 363
rect 917 317 963 363
rect 1037 317 1083 363
rect 1157 317 1203 363
rect 1277 317 1323 363
rect 1397 317 1443 363
rect 1517 317 1563 363
rect 1637 317 1683 363
rect 1757 317 1803 363
rect 1877 317 1923 363
rect 77 197 123 243
rect 197 197 243 243
rect 317 197 363 243
rect 437 197 483 243
rect 557 197 603 243
rect 677 197 723 243
rect 797 197 843 243
rect 917 197 963 243
rect 1037 197 1083 243
rect 1157 197 1203 243
rect 1277 197 1323 243
rect 1397 197 1443 243
rect 1517 197 1563 243
rect 1637 197 1683 243
rect 1757 197 1803 243
rect 1877 197 1923 243
rect 77 77 123 123
rect 197 77 243 123
rect 317 77 363 123
rect 437 77 483 123
rect 557 77 603 123
rect 677 77 723 123
rect 797 77 843 123
rect 917 77 963 123
rect 1037 77 1083 123
rect 1157 77 1203 123
rect 1277 77 1323 123
rect 1397 77 1443 123
rect 1517 77 1563 123
rect 1637 77 1683 123
rect 1757 77 1803 123
rect 1877 77 1923 123
<< psubdiff >>
rect -1264 3245 3264 3264
rect -1264 3199 -1091 3245
rect 3091 3199 3264 3245
rect -1264 3180 3264 3199
rect -1264 3091 -1180 3180
rect -1264 -1091 -1245 3091
rect -1199 -1091 -1180 3091
rect 3180 3091 3264 3180
rect -148 2129 2148 2148
rect -148 2083 -57 2129
rect 2057 2083 2148 2129
rect -148 2064 2148 2083
rect -148 2010 -64 2064
rect -148 -10 -129 2010
rect -83 -10 -64 2010
rect 2064 2010 2148 2064
rect -148 -64 -64 -10
rect 2064 -10 2083 2010
rect 2129 -10 2148 2010
rect 2064 -64 2148 -10
rect -148 -148 2148 -64
rect -1264 -1180 -1180 -1091
rect 3180 -1091 3199 3091
rect 3245 -1091 3264 3091
rect 3180 -1180 3264 -1091
rect -1264 -1199 3264 -1180
rect -1264 -1245 -1091 -1199
rect -763 -1245 2763 -1199
rect 3091 -1245 3264 -1199
rect -1264 -1264 3264 -1245
<< nsubdiff >>
rect -296 2277 2296 2296
rect -296 2231 -151 2277
rect 2151 2231 2296 2277
rect -296 2212 2296 2231
rect -296 2198 -212 2212
rect -296 -198 -277 2198
rect -231 -198 -212 2198
rect 2212 2198 2296 2212
rect -296 -212 -212 -198
rect 2212 -198 2231 2198
rect 2277 -198 2296 2198
rect 2212 -212 2296 -198
rect -296 -296 2296 -212
<< psubdiffcont >>
rect -1091 3199 3091 3245
rect -1245 -1091 -1199 3091
rect -57 2083 2057 2129
rect -129 -10 -83 2010
rect 2083 -10 2129 2010
rect 3199 -1091 3245 3091
rect -1091 -1245 -763 -1199
rect 2763 -1245 3091 -1199
<< nsubdiffcont >>
rect -151 2231 2151 2277
rect -277 -198 -231 2198
rect 2231 -198 2277 2198
<< metal1 >>
rect -1264 3245 3264 3264
rect -1264 3199 -1091 3245
rect 3091 3199 3264 3245
rect -1264 3180 3264 3199
rect -1264 3091 -1180 3180
rect -1264 -1091 -1245 3091
rect -1199 -1091 -1180 3091
rect 3180 3091 3264 3180
rect -296 2277 2296 2296
rect -296 2231 -151 2277
rect 2151 2231 2296 2277
rect -296 2212 2296 2231
rect -296 2198 -212 2212
rect -296 -198 -277 2198
rect -231 -198 -212 2198
rect 2212 2198 2296 2212
rect -148 2129 2148 2148
rect -148 2083 -57 2129
rect 2057 2083 2148 2129
rect -148 2064 2148 2083
rect -148 2010 -64 2064
rect -148 -10 -129 2010
rect -83 -10 -64 2010
rect 2064 2010 2148 2064
rect 0 1923 2000 2000
rect 0 1877 77 1923
rect 123 1877 197 1923
rect 243 1877 317 1923
rect 363 1877 437 1923
rect 483 1877 557 1923
rect 603 1877 677 1923
rect 723 1877 797 1923
rect 843 1877 917 1923
rect 963 1877 1037 1923
rect 1083 1877 1157 1923
rect 1203 1877 1277 1923
rect 1323 1877 1397 1923
rect 1443 1877 1517 1923
rect 1563 1877 1637 1923
rect 1683 1877 1757 1923
rect 1803 1877 1877 1923
rect 1923 1877 2000 1923
rect 0 1803 2000 1877
rect 0 1757 77 1803
rect 123 1757 197 1803
rect 243 1757 317 1803
rect 363 1757 437 1803
rect 483 1757 557 1803
rect 603 1757 677 1803
rect 723 1757 797 1803
rect 843 1757 917 1803
rect 963 1757 1037 1803
rect 1083 1757 1157 1803
rect 1203 1757 1277 1803
rect 1323 1757 1397 1803
rect 1443 1757 1517 1803
rect 1563 1757 1637 1803
rect 1683 1757 1757 1803
rect 1803 1757 1877 1803
rect 1923 1757 2000 1803
rect 0 1683 2000 1757
rect 0 1637 77 1683
rect 123 1637 197 1683
rect 243 1637 317 1683
rect 363 1637 437 1683
rect 483 1637 557 1683
rect 603 1637 677 1683
rect 723 1637 797 1683
rect 843 1637 917 1683
rect 963 1637 1037 1683
rect 1083 1637 1157 1683
rect 1203 1637 1277 1683
rect 1323 1637 1397 1683
rect 1443 1637 1517 1683
rect 1563 1637 1637 1683
rect 1683 1637 1757 1683
rect 1803 1637 1877 1683
rect 1923 1637 2000 1683
rect 0 1563 2000 1637
rect 0 1517 77 1563
rect 123 1517 197 1563
rect 243 1517 317 1563
rect 363 1517 437 1563
rect 483 1517 557 1563
rect 603 1517 677 1563
rect 723 1517 797 1563
rect 843 1517 917 1563
rect 963 1517 1037 1563
rect 1083 1517 1157 1563
rect 1203 1517 1277 1563
rect 1323 1517 1397 1563
rect 1443 1517 1517 1563
rect 1563 1517 1637 1563
rect 1683 1517 1757 1563
rect 1803 1517 1877 1563
rect 1923 1517 2000 1563
rect 0 1443 2000 1517
rect 0 1397 77 1443
rect 123 1397 197 1443
rect 243 1397 317 1443
rect 363 1397 437 1443
rect 483 1397 557 1443
rect 603 1397 677 1443
rect 723 1397 797 1443
rect 843 1397 917 1443
rect 963 1397 1037 1443
rect 1083 1397 1157 1443
rect 1203 1397 1277 1443
rect 1323 1397 1397 1443
rect 1443 1397 1517 1443
rect 1563 1397 1637 1443
rect 1683 1397 1757 1443
rect 1803 1397 1877 1443
rect 1923 1397 2000 1443
rect 0 1323 2000 1397
rect 0 1277 77 1323
rect 123 1277 197 1323
rect 243 1277 317 1323
rect 363 1277 437 1323
rect 483 1277 557 1323
rect 603 1277 677 1323
rect 723 1277 797 1323
rect 843 1277 917 1323
rect 963 1277 1037 1323
rect 1083 1277 1157 1323
rect 1203 1277 1277 1323
rect 1323 1277 1397 1323
rect 1443 1277 1517 1323
rect 1563 1277 1637 1323
rect 1683 1277 1757 1323
rect 1803 1277 1877 1323
rect 1923 1277 2000 1323
rect 0 1203 2000 1277
rect 0 1157 77 1203
rect 123 1157 197 1203
rect 243 1157 317 1203
rect 363 1157 437 1203
rect 483 1157 557 1203
rect 603 1157 677 1203
rect 723 1157 797 1203
rect 843 1157 917 1203
rect 963 1157 1037 1203
rect 1083 1157 1157 1203
rect 1203 1157 1277 1203
rect 1323 1157 1397 1203
rect 1443 1157 1517 1203
rect 1563 1157 1637 1203
rect 1683 1157 1757 1203
rect 1803 1157 1877 1203
rect 1923 1157 2000 1203
rect 0 1083 2000 1157
rect 0 1037 77 1083
rect 123 1037 197 1083
rect 243 1037 317 1083
rect 363 1037 437 1083
rect 483 1037 557 1083
rect 603 1037 677 1083
rect 723 1037 797 1083
rect 843 1037 917 1083
rect 963 1037 1037 1083
rect 1083 1037 1157 1083
rect 1203 1037 1277 1083
rect 1323 1037 1397 1083
rect 1443 1037 1517 1083
rect 1563 1037 1637 1083
rect 1683 1037 1757 1083
rect 1803 1037 1877 1083
rect 1923 1037 2000 1083
rect 0 963 2000 1037
rect 0 917 77 963
rect 123 917 197 963
rect 243 917 317 963
rect 363 917 437 963
rect 483 917 557 963
rect 603 917 677 963
rect 723 917 797 963
rect 843 917 917 963
rect 963 917 1037 963
rect 1083 917 1157 963
rect 1203 917 1277 963
rect 1323 917 1397 963
rect 1443 917 1517 963
rect 1563 917 1637 963
rect 1683 917 1757 963
rect 1803 917 1877 963
rect 1923 917 2000 963
rect 0 843 2000 917
rect 0 797 77 843
rect 123 797 197 843
rect 243 797 317 843
rect 363 797 437 843
rect 483 797 557 843
rect 603 797 677 843
rect 723 797 797 843
rect 843 797 917 843
rect 963 797 1037 843
rect 1083 797 1157 843
rect 1203 797 1277 843
rect 1323 797 1397 843
rect 1443 797 1517 843
rect 1563 797 1637 843
rect 1683 797 1757 843
rect 1803 797 1877 843
rect 1923 797 2000 843
rect 0 723 2000 797
rect 0 677 77 723
rect 123 677 197 723
rect 243 677 317 723
rect 363 677 437 723
rect 483 677 557 723
rect 603 677 677 723
rect 723 677 797 723
rect 843 677 917 723
rect 963 677 1037 723
rect 1083 677 1157 723
rect 1203 677 1277 723
rect 1323 677 1397 723
rect 1443 677 1517 723
rect 1563 677 1637 723
rect 1683 677 1757 723
rect 1803 677 1877 723
rect 1923 677 2000 723
rect 0 603 2000 677
rect 0 557 77 603
rect 123 557 197 603
rect 243 557 317 603
rect 363 557 437 603
rect 483 557 557 603
rect 603 557 677 603
rect 723 557 797 603
rect 843 557 917 603
rect 963 557 1037 603
rect 1083 557 1157 603
rect 1203 557 1277 603
rect 1323 557 1397 603
rect 1443 557 1517 603
rect 1563 557 1637 603
rect 1683 557 1757 603
rect 1803 557 1877 603
rect 1923 557 2000 603
rect 0 483 2000 557
rect 0 437 77 483
rect 123 437 197 483
rect 243 437 317 483
rect 363 437 437 483
rect 483 437 557 483
rect 603 437 677 483
rect 723 437 797 483
rect 843 437 917 483
rect 963 437 1037 483
rect 1083 437 1157 483
rect 1203 437 1277 483
rect 1323 437 1397 483
rect 1443 437 1517 483
rect 1563 437 1637 483
rect 1683 437 1757 483
rect 1803 437 1877 483
rect 1923 437 2000 483
rect 0 363 2000 437
rect 0 317 77 363
rect 123 317 197 363
rect 243 317 317 363
rect 363 317 437 363
rect 483 317 557 363
rect 603 317 677 363
rect 723 317 797 363
rect 843 317 917 363
rect 963 317 1037 363
rect 1083 317 1157 363
rect 1203 317 1277 363
rect 1323 317 1397 363
rect 1443 317 1517 363
rect 1563 317 1637 363
rect 1683 317 1757 363
rect 1803 317 1877 363
rect 1923 317 2000 363
rect 0 243 2000 317
rect 0 197 77 243
rect 123 197 197 243
rect 243 197 317 243
rect 363 197 437 243
rect 483 197 557 243
rect 603 197 677 243
rect 723 197 797 243
rect 843 197 917 243
rect 963 197 1037 243
rect 1083 197 1157 243
rect 1203 197 1277 243
rect 1323 197 1397 243
rect 1443 197 1517 243
rect 1563 197 1637 243
rect 1683 197 1757 243
rect 1803 197 1877 243
rect 1923 197 2000 243
rect 0 123 2000 197
rect 0 77 77 123
rect 123 77 197 123
rect 243 77 317 123
rect 363 77 437 123
rect 483 77 557 123
rect 603 77 677 123
rect 723 77 797 123
rect 843 77 917 123
rect 963 77 1037 123
rect 1083 77 1157 123
rect 1203 77 1277 123
rect 1323 77 1397 123
rect 1443 77 1517 123
rect 1563 77 1637 123
rect 1683 77 1757 123
rect 1803 77 1877 123
rect 1923 77 2000 123
rect 0 0 2000 77
rect -148 -148 -64 -10
rect 2064 -10 2083 2010
rect 2129 -10 2148 2010
rect 2064 -148 2148 -10
rect -296 -296 -212 -198
rect 2212 -198 2231 2198
rect 2277 -198 2296 2198
rect 2212 -296 2296 -198
rect -1264 -1180 -1180 -1091
rect 3180 -1091 3199 3091
rect 3245 -1091 3264 3091
rect 3180 -1180 3264 -1091
rect -1264 -1199 -680 -1180
rect -1264 -1245 -1091 -1199
rect -763 -1245 -680 -1199
rect -1264 -1264 -680 -1245
rect 2680 -1199 3264 -1180
rect 2680 -1245 2763 -1199
rect 3091 -1245 3264 -1199
rect 2680 -1264 3264 -1245
<< labels >>
flabel metal1 1001 999 1001 999 0 FreeSans 400 0 0 0 E
flabel metal1 -103 -97 -103 -97 0 FreeSans 400 0 0 0 B
flabel metal1 2105 -99 2105 -99 0 FreeSans 400 0 0 0 B
flabel metal1 2110 2108 2110 2108 0 FreeSans 400 0 0 0 B
flabel metal1 -251 2252 -251 2252 0 FreeSans 400 0 0 0 C
flabel metal1 2254 -247 2254 -247 0 FreeSans 400 0 0 0 C
flabel metal1 2257 2257 2257 2257 0 FreeSans 400 0 0 0 C
flabel metal1 3221 3221 3221 3221 0 FreeSans 400 0 0 0 S
flabel metal1 3214 -1219 3214 -1219 0 FreeSans 400 0 0 0 S
flabel metal1 3214 -1219 3214 -1219 0 FreeSans 400 0 0 0 S
flabel metal1 -1219 -1211 -1219 -1211 0 FreeSans 400 0 0 0 S
flabel metal1 -1219 -1211 -1219 -1211 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 37868
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_10p00x10p00.gds
string GDS_START 112
string gencell npn_10p00x10p00
string library gf180mcu
string parameter m=1
<< end >>
