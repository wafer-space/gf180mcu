magic
tech gf180mcuD
timestamp 1755724134
<< properties >>
string GDS_END 1061838
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1059594
<< end >>
