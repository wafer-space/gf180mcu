magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 7254 1094
<< pwell >>
rect -86 -86 7254 453
<< mvnmos >>
rect 124 69 324 333
rect 572 69 772 333
rect 1020 69 1220 333
rect 1468 69 1668 333
rect 1916 69 2116 333
rect 2364 69 2564 333
rect 2812 69 3012 333
rect 3260 69 3460 333
rect 3708 69 3908 333
rect 4156 69 4356 333
rect 4604 69 4804 333
rect 5052 69 5252 333
rect 5500 69 5700 333
rect 5948 69 6148 333
rect 6396 69 6596 333
rect 6844 69 7044 333
<< mvpmos >>
rect 124 573 324 939
rect 572 573 772 939
rect 1020 573 1220 939
rect 1468 573 1668 939
rect 1916 573 2116 939
rect 2364 573 2564 939
rect 2812 573 3012 939
rect 3260 573 3460 939
rect 3708 573 3908 939
rect 4156 573 4356 939
rect 4604 573 4804 939
rect 5052 573 5252 939
rect 5500 573 5700 939
rect 5948 573 6148 939
rect 6396 573 6596 939
rect 6844 573 7044 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 324 287 412 333
rect 324 147 353 287
rect 399 147 412 287
rect 324 69 412 147
rect 484 287 572 333
rect 484 147 497 287
rect 543 147 572 287
rect 484 69 572 147
rect 772 287 860 333
rect 772 147 801 287
rect 847 147 860 287
rect 772 69 860 147
rect 932 287 1020 333
rect 932 147 945 287
rect 991 147 1020 287
rect 932 69 1020 147
rect 1220 287 1308 333
rect 1220 147 1249 287
rect 1295 147 1308 287
rect 1220 69 1308 147
rect 1380 287 1468 333
rect 1380 147 1393 287
rect 1439 147 1468 287
rect 1380 69 1468 147
rect 1668 287 1756 333
rect 1668 147 1697 287
rect 1743 147 1756 287
rect 1668 69 1756 147
rect 1828 287 1916 333
rect 1828 147 1841 287
rect 1887 147 1916 287
rect 1828 69 1916 147
rect 2116 287 2204 333
rect 2116 147 2145 287
rect 2191 147 2204 287
rect 2116 69 2204 147
rect 2276 287 2364 333
rect 2276 147 2289 287
rect 2335 147 2364 287
rect 2276 69 2364 147
rect 2564 287 2652 333
rect 2564 147 2593 287
rect 2639 147 2652 287
rect 2564 69 2652 147
rect 2724 287 2812 333
rect 2724 147 2737 287
rect 2783 147 2812 287
rect 2724 69 2812 147
rect 3012 287 3100 333
rect 3012 147 3041 287
rect 3087 147 3100 287
rect 3012 69 3100 147
rect 3172 287 3260 333
rect 3172 147 3185 287
rect 3231 147 3260 287
rect 3172 69 3260 147
rect 3460 287 3548 333
rect 3460 147 3489 287
rect 3535 147 3548 287
rect 3460 69 3548 147
rect 3620 287 3708 333
rect 3620 147 3633 287
rect 3679 147 3708 287
rect 3620 69 3708 147
rect 3908 287 3996 333
rect 3908 147 3937 287
rect 3983 147 3996 287
rect 3908 69 3996 147
rect 4068 287 4156 333
rect 4068 147 4081 287
rect 4127 147 4156 287
rect 4068 69 4156 147
rect 4356 287 4444 333
rect 4356 147 4385 287
rect 4431 147 4444 287
rect 4356 69 4444 147
rect 4516 287 4604 333
rect 4516 147 4529 287
rect 4575 147 4604 287
rect 4516 69 4604 147
rect 4804 287 4892 333
rect 4804 147 4833 287
rect 4879 147 4892 287
rect 4804 69 4892 147
rect 4964 287 5052 333
rect 4964 147 4977 287
rect 5023 147 5052 287
rect 4964 69 5052 147
rect 5252 287 5340 333
rect 5252 147 5281 287
rect 5327 147 5340 287
rect 5252 69 5340 147
rect 5412 287 5500 333
rect 5412 147 5425 287
rect 5471 147 5500 287
rect 5412 69 5500 147
rect 5700 287 5788 333
rect 5700 147 5729 287
rect 5775 147 5788 287
rect 5700 69 5788 147
rect 5860 287 5948 333
rect 5860 147 5873 287
rect 5919 147 5948 287
rect 5860 69 5948 147
rect 6148 287 6236 333
rect 6148 147 6177 287
rect 6223 147 6236 287
rect 6148 69 6236 147
rect 6308 287 6396 333
rect 6308 147 6321 287
rect 6367 147 6396 287
rect 6308 69 6396 147
rect 6596 287 6684 333
rect 6596 147 6625 287
rect 6671 147 6684 287
rect 6596 69 6684 147
rect 6756 287 6844 333
rect 6756 147 6769 287
rect 6815 147 6844 287
rect 6756 69 6844 147
rect 7044 287 7132 333
rect 7044 147 7073 287
rect 7119 147 7132 287
rect 7044 69 7132 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 324 861 412 939
rect 324 721 353 861
rect 399 721 412 861
rect 324 573 412 721
rect 484 861 572 939
rect 484 721 497 861
rect 543 721 572 861
rect 484 573 572 721
rect 772 861 860 939
rect 772 721 801 861
rect 847 721 860 861
rect 772 573 860 721
rect 932 861 1020 939
rect 932 721 945 861
rect 991 721 1020 861
rect 932 573 1020 721
rect 1220 861 1308 939
rect 1220 721 1249 861
rect 1295 721 1308 861
rect 1220 573 1308 721
rect 1380 861 1468 939
rect 1380 721 1393 861
rect 1439 721 1468 861
rect 1380 573 1468 721
rect 1668 861 1756 939
rect 1668 721 1697 861
rect 1743 721 1756 861
rect 1668 573 1756 721
rect 1828 861 1916 939
rect 1828 721 1841 861
rect 1887 721 1916 861
rect 1828 573 1916 721
rect 2116 861 2204 939
rect 2116 721 2145 861
rect 2191 721 2204 861
rect 2116 573 2204 721
rect 2276 861 2364 939
rect 2276 721 2289 861
rect 2335 721 2364 861
rect 2276 573 2364 721
rect 2564 861 2652 939
rect 2564 721 2593 861
rect 2639 721 2652 861
rect 2564 573 2652 721
rect 2724 861 2812 939
rect 2724 721 2737 861
rect 2783 721 2812 861
rect 2724 573 2812 721
rect 3012 861 3100 939
rect 3012 721 3041 861
rect 3087 721 3100 861
rect 3012 573 3100 721
rect 3172 861 3260 939
rect 3172 721 3185 861
rect 3231 721 3260 861
rect 3172 573 3260 721
rect 3460 861 3548 939
rect 3460 721 3489 861
rect 3535 721 3548 861
rect 3460 573 3548 721
rect 3620 861 3708 939
rect 3620 721 3633 861
rect 3679 721 3708 861
rect 3620 573 3708 721
rect 3908 861 3996 939
rect 3908 721 3937 861
rect 3983 721 3996 861
rect 3908 573 3996 721
rect 4068 861 4156 939
rect 4068 721 4081 861
rect 4127 721 4156 861
rect 4068 573 4156 721
rect 4356 861 4444 939
rect 4356 721 4385 861
rect 4431 721 4444 861
rect 4356 573 4444 721
rect 4516 861 4604 939
rect 4516 721 4529 861
rect 4575 721 4604 861
rect 4516 573 4604 721
rect 4804 861 4892 939
rect 4804 721 4833 861
rect 4879 721 4892 861
rect 4804 573 4892 721
rect 4964 861 5052 939
rect 4964 721 4977 861
rect 5023 721 5052 861
rect 4964 573 5052 721
rect 5252 861 5340 939
rect 5252 721 5281 861
rect 5327 721 5340 861
rect 5252 573 5340 721
rect 5412 861 5500 939
rect 5412 721 5425 861
rect 5471 721 5500 861
rect 5412 573 5500 721
rect 5700 861 5788 939
rect 5700 721 5729 861
rect 5775 721 5788 861
rect 5700 573 5788 721
rect 5860 861 5948 939
rect 5860 721 5873 861
rect 5919 721 5948 861
rect 5860 573 5948 721
rect 6148 861 6236 939
rect 6148 721 6177 861
rect 6223 721 6236 861
rect 6148 573 6236 721
rect 6308 861 6396 939
rect 6308 721 6321 861
rect 6367 721 6396 861
rect 6308 573 6396 721
rect 6596 861 6684 939
rect 6596 721 6625 861
rect 6671 721 6684 861
rect 6596 573 6684 721
rect 6756 861 6844 939
rect 6756 721 6769 861
rect 6815 721 6844 861
rect 6756 573 6844 721
rect 7044 861 7132 939
rect 7044 721 7073 861
rect 7119 721 7132 861
rect 7044 573 7132 721
<< mvndiffc >>
rect 49 147 95 287
rect 353 147 399 287
rect 497 147 543 287
rect 801 147 847 287
rect 945 147 991 287
rect 1249 147 1295 287
rect 1393 147 1439 287
rect 1697 147 1743 287
rect 1841 147 1887 287
rect 2145 147 2191 287
rect 2289 147 2335 287
rect 2593 147 2639 287
rect 2737 147 2783 287
rect 3041 147 3087 287
rect 3185 147 3231 287
rect 3489 147 3535 287
rect 3633 147 3679 287
rect 3937 147 3983 287
rect 4081 147 4127 287
rect 4385 147 4431 287
rect 4529 147 4575 287
rect 4833 147 4879 287
rect 4977 147 5023 287
rect 5281 147 5327 287
rect 5425 147 5471 287
rect 5729 147 5775 287
rect 5873 147 5919 287
rect 6177 147 6223 287
rect 6321 147 6367 287
rect 6625 147 6671 287
rect 6769 147 6815 287
rect 7073 147 7119 287
<< mvpdiffc >>
rect 49 721 95 861
rect 353 721 399 861
rect 497 721 543 861
rect 801 721 847 861
rect 945 721 991 861
rect 1249 721 1295 861
rect 1393 721 1439 861
rect 1697 721 1743 861
rect 1841 721 1887 861
rect 2145 721 2191 861
rect 2289 721 2335 861
rect 2593 721 2639 861
rect 2737 721 2783 861
rect 3041 721 3087 861
rect 3185 721 3231 861
rect 3489 721 3535 861
rect 3633 721 3679 861
rect 3937 721 3983 861
rect 4081 721 4127 861
rect 4385 721 4431 861
rect 4529 721 4575 861
rect 4833 721 4879 861
rect 4977 721 5023 861
rect 5281 721 5327 861
rect 5425 721 5471 861
rect 5729 721 5775 861
rect 5873 721 5919 861
rect 6177 721 6223 861
rect 6321 721 6367 861
rect 6625 721 6671 861
rect 6769 721 6815 861
rect 7073 721 7119 861
<< polysilicon >>
rect 124 939 324 983
rect 572 939 772 983
rect 1020 939 1220 983
rect 1468 939 1668 983
rect 1916 939 2116 983
rect 2364 939 2564 983
rect 2812 939 3012 983
rect 3260 939 3460 983
rect 3708 939 3908 983
rect 4156 939 4356 983
rect 4604 939 4804 983
rect 5052 939 5252 983
rect 5500 939 5700 983
rect 5948 939 6148 983
rect 6396 939 6596 983
rect 6844 939 7044 983
rect 124 540 324 573
rect 124 494 265 540
rect 311 494 324 540
rect 124 481 324 494
rect 572 540 772 573
rect 572 494 713 540
rect 759 494 772 540
rect 572 481 772 494
rect 1020 540 1220 573
rect 1020 494 1161 540
rect 1207 494 1220 540
rect 1020 481 1220 494
rect 1468 540 1668 573
rect 1468 494 1609 540
rect 1655 494 1668 540
rect 1468 481 1668 494
rect 1916 540 2116 573
rect 1916 494 2057 540
rect 2103 494 2116 540
rect 1916 481 2116 494
rect 2364 540 2564 573
rect 2364 494 2505 540
rect 2551 494 2564 540
rect 2364 481 2564 494
rect 2812 540 3012 573
rect 2812 494 2953 540
rect 2999 494 3012 540
rect 2812 481 3012 494
rect 3260 540 3460 573
rect 3260 494 3401 540
rect 3447 494 3460 540
rect 3260 481 3460 494
rect 3708 540 3908 573
rect 3708 494 3849 540
rect 3895 494 3908 540
rect 3708 481 3908 494
rect 4156 540 4356 573
rect 4156 494 4297 540
rect 4343 494 4356 540
rect 4156 481 4356 494
rect 4604 540 4804 573
rect 4604 494 4745 540
rect 4791 494 4804 540
rect 4604 481 4804 494
rect 5052 540 5252 573
rect 5052 494 5193 540
rect 5239 494 5252 540
rect 5052 481 5252 494
rect 5500 540 5700 573
rect 5500 494 5641 540
rect 5687 494 5700 540
rect 5500 481 5700 494
rect 5948 540 6148 573
rect 5948 494 6089 540
rect 6135 494 6148 540
rect 5948 481 6148 494
rect 6396 540 6596 573
rect 6396 494 6537 540
rect 6583 494 6596 540
rect 6396 481 6596 494
rect 6844 540 7044 573
rect 6844 494 6985 540
rect 7031 494 7044 540
rect 6844 481 7044 494
rect 124 412 324 425
rect 124 366 137 412
rect 183 366 324 412
rect 124 333 324 366
rect 572 412 772 425
rect 572 366 585 412
rect 631 366 772 412
rect 572 333 772 366
rect 1020 412 1220 425
rect 1020 366 1033 412
rect 1079 366 1220 412
rect 1020 333 1220 366
rect 1468 412 1668 425
rect 1468 366 1481 412
rect 1527 366 1668 412
rect 1468 333 1668 366
rect 1916 412 2116 425
rect 1916 366 1929 412
rect 1975 366 2116 412
rect 1916 333 2116 366
rect 2364 412 2564 425
rect 2364 366 2377 412
rect 2423 366 2564 412
rect 2364 333 2564 366
rect 2812 412 3012 425
rect 2812 366 2825 412
rect 2871 366 3012 412
rect 2812 333 3012 366
rect 3260 412 3460 425
rect 3260 366 3273 412
rect 3319 366 3460 412
rect 3260 333 3460 366
rect 3708 412 3908 425
rect 3708 366 3721 412
rect 3767 366 3908 412
rect 3708 333 3908 366
rect 4156 412 4356 425
rect 4156 366 4169 412
rect 4215 366 4356 412
rect 4156 333 4356 366
rect 4604 412 4804 425
rect 4604 366 4617 412
rect 4663 366 4804 412
rect 4604 333 4804 366
rect 5052 412 5252 425
rect 5052 366 5065 412
rect 5111 366 5252 412
rect 5052 333 5252 366
rect 5500 412 5700 425
rect 5500 366 5513 412
rect 5559 366 5700 412
rect 5500 333 5700 366
rect 5948 412 6148 425
rect 5948 366 5961 412
rect 6007 366 6148 412
rect 5948 333 6148 366
rect 6396 412 6596 425
rect 6396 366 6409 412
rect 6455 366 6596 412
rect 6396 333 6596 366
rect 6844 412 7044 425
rect 6844 366 6857 412
rect 6903 366 7044 412
rect 6844 333 7044 366
rect 124 25 324 69
rect 572 25 772 69
rect 1020 25 1220 69
rect 1468 25 1668 69
rect 1916 25 2116 69
rect 2364 25 2564 69
rect 2812 25 3012 69
rect 3260 25 3460 69
rect 3708 25 3908 69
rect 4156 25 4356 69
rect 4604 25 4804 69
rect 5052 25 5252 69
rect 5500 25 5700 69
rect 5948 25 6148 69
rect 6396 25 6596 69
rect 6844 25 7044 69
<< polycontact >>
rect 265 494 311 540
rect 713 494 759 540
rect 1161 494 1207 540
rect 1609 494 1655 540
rect 2057 494 2103 540
rect 2505 494 2551 540
rect 2953 494 2999 540
rect 3401 494 3447 540
rect 3849 494 3895 540
rect 4297 494 4343 540
rect 4745 494 4791 540
rect 5193 494 5239 540
rect 5641 494 5687 540
rect 6089 494 6135 540
rect 6537 494 6583 540
rect 6985 494 7031 540
rect 137 366 183 412
rect 585 366 631 412
rect 1033 366 1079 412
rect 1481 366 1527 412
rect 1929 366 1975 412
rect 2377 366 2423 412
rect 2825 366 2871 412
rect 3273 366 3319 412
rect 3721 366 3767 412
rect 4169 366 4215 412
rect 4617 366 4663 412
rect 5065 366 5111 412
rect 5513 366 5559 412
rect 5961 366 6007 412
rect 6409 366 6455 412
rect 6857 366 6903 412
<< metal1 >>
rect 0 918 7168 1098
rect 49 861 95 872
rect 49 412 95 721
rect 353 861 399 918
rect 353 710 399 721
rect 497 861 543 872
rect 265 540 311 551
rect 49 366 137 412
rect 183 366 194 412
rect 265 298 311 494
rect 497 412 543 721
rect 801 861 847 918
rect 801 710 847 721
rect 945 861 991 872
rect 713 540 759 551
rect 497 366 585 412
rect 631 366 642 412
rect 713 298 759 494
rect 945 412 991 721
rect 1249 861 1295 918
rect 1249 710 1295 721
rect 1393 861 1439 872
rect 1161 540 1207 551
rect 945 366 1033 412
rect 1079 366 1090 412
rect 1161 298 1207 494
rect 1393 412 1439 721
rect 1697 861 1743 918
rect 1697 710 1743 721
rect 1841 861 1887 872
rect 1609 540 1655 551
rect 1393 366 1481 412
rect 1527 366 1538 412
rect 1609 298 1655 494
rect 1841 412 1887 721
rect 2145 861 2191 918
rect 2145 710 2191 721
rect 2289 861 2335 872
rect 2057 540 2103 551
rect 1841 366 1929 412
rect 1975 366 1986 412
rect 2057 298 2103 494
rect 2289 412 2335 721
rect 2593 861 2639 918
rect 2593 710 2639 721
rect 2737 861 2783 872
rect 2505 540 2551 551
rect 2289 366 2377 412
rect 2423 366 2434 412
rect 2505 298 2551 494
rect 2737 412 2783 721
rect 3041 861 3087 918
rect 3041 710 3087 721
rect 3185 861 3231 872
rect 2953 540 2999 551
rect 2737 366 2825 412
rect 2871 366 2882 412
rect 2953 298 2999 494
rect 3185 412 3231 721
rect 3489 861 3535 918
rect 3489 710 3535 721
rect 3633 861 3679 872
rect 3401 540 3447 551
rect 3185 366 3273 412
rect 3319 366 3330 412
rect 3401 298 3447 494
rect 3633 412 3679 721
rect 3937 861 3983 918
rect 3937 710 3983 721
rect 4081 861 4127 872
rect 3849 540 3895 551
rect 3633 366 3721 412
rect 3767 366 3778 412
rect 3849 298 3895 494
rect 4081 412 4127 721
rect 4385 861 4431 918
rect 4385 710 4431 721
rect 4529 861 4575 872
rect 4297 540 4343 551
rect 4081 366 4169 412
rect 4215 366 4226 412
rect 4297 298 4343 494
rect 4529 412 4575 721
rect 4833 861 4879 918
rect 4833 710 4879 721
rect 4977 861 5023 872
rect 4745 540 4791 551
rect 4529 366 4617 412
rect 4663 366 4674 412
rect 4745 298 4791 494
rect 4977 412 5023 721
rect 5281 861 5327 918
rect 5281 710 5327 721
rect 5425 861 5471 872
rect 5193 540 5239 551
rect 4977 366 5065 412
rect 5111 366 5122 412
rect 5193 298 5239 494
rect 5425 412 5471 721
rect 5729 861 5775 918
rect 5729 710 5775 721
rect 5873 861 5919 872
rect 5641 540 5687 551
rect 5425 366 5513 412
rect 5559 366 5570 412
rect 5641 298 5687 494
rect 5873 412 5919 721
rect 6177 861 6223 918
rect 6177 710 6223 721
rect 6321 861 6367 872
rect 6089 540 6135 551
rect 5873 366 5961 412
rect 6007 366 6018 412
rect 6089 298 6135 494
rect 6321 412 6367 721
rect 6625 861 6671 918
rect 6625 710 6671 721
rect 6769 861 6815 872
rect 6537 540 6583 551
rect 6321 366 6409 412
rect 6455 366 6466 412
rect 6537 298 6583 494
rect 6769 412 6815 721
rect 7073 861 7119 918
rect 7073 710 7119 721
rect 6985 540 7031 551
rect 6769 366 6857 412
rect 6903 366 6914 412
rect 6985 298 7031 494
rect 49 287 95 298
rect 265 287 399 298
rect 265 252 353 287
rect 49 90 95 147
rect 353 136 399 147
rect 497 287 543 298
rect 713 287 847 298
rect 713 252 801 287
rect 497 90 543 147
rect 801 136 847 147
rect 945 287 991 298
rect 1161 287 1295 298
rect 1161 252 1249 287
rect 945 90 991 147
rect 1249 136 1295 147
rect 1393 287 1439 298
rect 1609 287 1743 298
rect 1609 252 1697 287
rect 1393 90 1439 147
rect 1697 136 1743 147
rect 1841 287 1887 298
rect 2057 287 2191 298
rect 2057 252 2145 287
rect 1841 90 1887 147
rect 2145 136 2191 147
rect 2289 287 2335 298
rect 2505 287 2639 298
rect 2505 252 2593 287
rect 2289 90 2335 147
rect 2593 136 2639 147
rect 2737 287 2783 298
rect 2953 287 3087 298
rect 2953 252 3041 287
rect 2737 90 2783 147
rect 3041 136 3087 147
rect 3185 287 3231 298
rect 3401 287 3535 298
rect 3401 252 3489 287
rect 3185 90 3231 147
rect 3489 136 3535 147
rect 3633 287 3679 298
rect 3849 287 3983 298
rect 3849 252 3937 287
rect 3633 90 3679 147
rect 3937 136 3983 147
rect 4081 287 4127 298
rect 4297 287 4431 298
rect 4297 252 4385 287
rect 4081 90 4127 147
rect 4385 136 4431 147
rect 4529 287 4575 298
rect 4745 287 4879 298
rect 4745 252 4833 287
rect 4529 90 4575 147
rect 4833 136 4879 147
rect 4977 287 5023 298
rect 5193 287 5327 298
rect 5193 252 5281 287
rect 4977 90 5023 147
rect 5281 136 5327 147
rect 5425 287 5471 298
rect 5641 287 5775 298
rect 5641 252 5729 287
rect 5425 90 5471 147
rect 5729 136 5775 147
rect 5873 287 5919 298
rect 6089 287 6223 298
rect 6089 252 6177 287
rect 5873 90 5919 147
rect 6177 136 6223 147
rect 6321 287 6367 298
rect 6537 287 6671 298
rect 6537 252 6625 287
rect 6321 90 6367 147
rect 6625 136 6671 147
rect 6769 287 6815 298
rect 6985 287 7119 298
rect 6985 252 7073 287
rect 6769 90 6815 147
rect 7073 136 7119 147
rect 0 -90 7168 90
<< labels >>
flabel metal1 s 0 918 7168 1098 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 6769 90 6815 298 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 7073 710 7119 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6625 710 6671 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6177 710 6223 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5729 710 5775 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5281 710 5327 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4833 710 4879 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4385 710 4431 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3937 710 3983 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3489 710 3535 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3041 710 3087 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2593 710 2639 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2145 710 2191 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 710 1743 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 710 1295 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 710 847 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 710 399 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6321 90 6367 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5873 90 5919 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5425 90 5471 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4977 90 5023 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 90 4575 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4081 90 4127 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3633 90 3679 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3185 90 3231 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2737 90 2783 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 7168 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 7168 1008
string GDS_END 814884
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 795546
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
