magic
tech gf180mcuD
timestamp 1755724134
<< properties >>
string GDS_END 11705116
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 11664664
<< end >>
