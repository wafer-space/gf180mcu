magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 377 4342 870
rect -86 352 1453 377
rect 4070 352 4342 377
<< pwell >>
rect 1453 352 4070 377
rect -86 -86 4342 352
<< mvnmos >>
rect 150 124 270 217
rect 374 124 494 217
rect 742 156 862 228
rect 966 156 1086 228
rect 1190 156 1310 228
rect 1358 156 1478 228
rect 1670 185 1790 257
rect 1894 185 2014 257
rect 2118 185 2238 257
rect 2432 68 2552 257
rect 2656 68 2776 257
rect 3116 68 3236 232
rect 3428 68 3548 232
rect 3652 68 3772 232
rect 3964 68 4084 232
<< mvpmos >>
rect 170 472 270 645
rect 374 472 474 645
rect 766 500 866 599
rect 970 500 1070 599
rect 1201 500 1301 599
rect 1378 500 1478 599
rect 1670 500 1770 599
rect 1893 500 1993 599
rect 2204 500 2304 599
rect 2452 500 2552 715
rect 2656 500 2756 715
rect 3136 497 3236 716
rect 3428 497 3528 716
rect 3632 497 3732 716
rect 3880 497 3980 716
<< mvndiff >>
rect 1538 228 1670 257
rect 62 204 150 217
rect 62 158 75 204
rect 121 158 150 204
rect 62 124 150 158
rect 270 183 374 217
rect 270 137 299 183
rect 345 137 374 183
rect 270 124 374 137
rect 494 204 582 217
rect 494 158 523 204
rect 569 158 582 204
rect 494 124 582 158
rect 654 215 742 228
rect 654 169 667 215
rect 713 169 742 215
rect 654 156 742 169
rect 862 215 966 228
rect 862 169 891 215
rect 937 169 966 215
rect 862 156 966 169
rect 1086 215 1190 228
rect 1086 169 1115 215
rect 1161 169 1190 215
rect 1086 156 1190 169
rect 1310 156 1358 228
rect 1478 185 1670 228
rect 1790 244 1894 257
rect 1790 198 1819 244
rect 1865 198 1894 244
rect 1790 185 1894 198
rect 2014 244 2118 257
rect 2014 198 2043 244
rect 2089 198 2118 244
rect 2014 185 2118 198
rect 2238 192 2432 257
rect 2238 185 2349 192
rect 1478 162 1610 185
rect 1478 156 1551 162
rect 1538 116 1551 156
rect 1597 116 1610 162
rect 1538 103 1610 116
rect 2336 146 2349 185
rect 2395 146 2432 192
rect 2336 68 2432 146
rect 2552 127 2656 257
rect 2552 81 2581 127
rect 2627 81 2656 127
rect 2552 68 2656 81
rect 2776 244 2900 257
rect 2776 198 2841 244
rect 2887 198 2900 244
rect 3296 244 3368 257
rect 3296 232 3309 244
rect 2776 68 2900 198
rect 3028 127 3116 232
rect 3028 81 3041 127
rect 3087 81 3116 127
rect 3028 68 3116 81
rect 3236 198 3309 232
rect 3355 232 3368 244
rect 3832 244 3904 257
rect 3832 232 3845 244
rect 3355 198 3428 232
rect 3236 68 3428 198
rect 3548 127 3652 232
rect 3548 81 3577 127
rect 3623 81 3652 127
rect 3548 68 3652 81
rect 3772 198 3845 232
rect 3891 232 3904 244
rect 3891 198 3964 232
rect 3772 68 3964 198
rect 4084 142 4172 232
rect 4084 96 4113 142
rect 4159 96 4172 142
rect 4084 68 4172 96
<< mvpdiff >>
rect 634 647 706 660
rect 82 632 170 645
rect 82 492 95 632
rect 141 492 170 632
rect 82 472 170 492
rect 270 632 374 645
rect 270 586 299 632
rect 345 586 374 632
rect 270 472 374 586
rect 474 632 562 645
rect 474 492 503 632
rect 549 492 562 632
rect 634 601 647 647
rect 693 601 706 647
rect 634 599 706 601
rect 2364 609 2452 715
rect 2364 599 2377 609
rect 634 500 766 599
rect 866 575 970 599
rect 866 529 895 575
rect 941 529 970 575
rect 866 500 970 529
rect 1070 559 1201 599
rect 1070 513 1126 559
rect 1172 513 1201 559
rect 1070 500 1201 513
rect 1301 500 1378 599
rect 1478 586 1670 599
rect 1478 540 1552 586
rect 1598 540 1670 586
rect 1478 500 1670 540
rect 1770 575 1893 599
rect 1770 529 1818 575
rect 1864 529 1893 575
rect 1770 500 1893 529
rect 1993 575 2204 599
rect 1993 529 2043 575
rect 2089 529 2204 575
rect 1993 500 2204 529
rect 2304 563 2377 599
rect 2423 563 2452 609
rect 2304 500 2452 563
rect 2552 702 2656 715
rect 2552 656 2581 702
rect 2627 656 2656 702
rect 2552 500 2656 656
rect 2756 559 2888 715
rect 2756 513 2829 559
rect 2875 513 2888 559
rect 2756 500 2888 513
rect 3048 703 3136 716
rect 3048 563 3061 703
rect 3107 563 3136 703
rect 474 472 562 492
rect 3048 497 3136 563
rect 3236 586 3428 716
rect 3236 540 3309 586
rect 3355 540 3428 586
rect 3236 497 3428 540
rect 3528 703 3632 716
rect 3528 657 3557 703
rect 3603 657 3632 703
rect 3528 497 3632 657
rect 3732 586 3880 716
rect 3732 540 3785 586
rect 3831 540 3880 586
rect 3732 497 3880 540
rect 3980 703 4172 716
rect 3980 563 4113 703
rect 4159 563 4172 703
rect 3980 497 4172 563
<< mvndiffc >>
rect 75 158 121 204
rect 299 137 345 183
rect 523 158 569 204
rect 667 169 713 215
rect 891 169 937 215
rect 1115 169 1161 215
rect 1819 198 1865 244
rect 2043 198 2089 244
rect 1551 116 1597 162
rect 2349 146 2395 192
rect 2581 81 2627 127
rect 2841 198 2887 244
rect 3041 81 3087 127
rect 3309 198 3355 244
rect 3577 81 3623 127
rect 3845 198 3891 244
rect 4113 96 4159 142
<< mvpdiffc >>
rect 95 492 141 632
rect 299 586 345 632
rect 503 492 549 632
rect 647 601 693 647
rect 895 529 941 575
rect 1126 513 1172 559
rect 1552 540 1598 586
rect 1818 529 1864 575
rect 2043 529 2089 575
rect 2377 563 2423 609
rect 2581 656 2627 702
rect 2829 513 2875 559
rect 3061 563 3107 703
rect 3309 540 3355 586
rect 3557 657 3603 703
rect 3785 540 3831 586
rect 4113 563 4159 703
<< polysilicon >>
rect 374 720 1070 760
rect 170 645 270 690
rect 374 645 474 720
rect 766 599 866 643
rect 970 599 1070 720
rect 1201 720 1993 760
rect 1201 678 1301 720
rect 1201 632 1214 678
rect 1260 632 1301 678
rect 1201 599 1301 632
rect 1378 599 1478 643
rect 1670 599 1770 643
rect 1893 599 1993 720
rect 2452 715 2552 760
rect 2656 715 2756 760
rect 3136 716 3236 760
rect 3428 716 3528 760
rect 3632 716 3732 760
rect 3880 716 3980 760
rect 2204 599 2304 643
rect 170 412 270 472
rect 170 366 183 412
rect 229 366 270 412
rect 170 261 270 366
rect 150 217 270 261
rect 374 326 474 472
rect 374 280 387 326
rect 433 280 474 326
rect 374 261 474 280
rect 766 415 866 500
rect 970 456 1070 500
rect 766 369 807 415
rect 853 369 866 415
rect 1201 408 1301 500
rect 766 288 866 369
rect 966 368 1301 408
rect 1378 467 1478 500
rect 1378 421 1419 467
rect 1465 421 1478 467
rect 766 272 862 288
rect 374 217 494 261
rect 742 228 862 272
rect 966 228 1086 368
rect 1190 307 1310 320
rect 1190 261 1218 307
rect 1264 261 1310 307
rect 1378 272 1478 421
rect 1190 228 1310 261
rect 1358 228 1478 272
rect 1670 346 1770 500
rect 1893 399 1993 500
rect 2204 456 2304 500
rect 2232 408 2304 456
rect 1893 359 2158 399
rect 1670 300 1683 346
rect 1729 301 1770 346
rect 2118 301 2158 359
rect 2232 362 2245 408
rect 2291 362 2304 408
rect 2232 349 2304 362
rect 2452 346 2552 500
rect 2452 301 2493 346
rect 1729 300 1790 301
rect 1670 257 1790 300
rect 1894 257 2014 301
rect 2118 257 2238 301
rect 2432 300 2493 301
rect 2539 300 2552 346
rect 2432 257 2552 300
rect 2656 467 2756 500
rect 2656 421 2697 467
rect 2743 421 2756 467
rect 2656 301 2756 421
rect 3136 416 3236 497
rect 3428 416 3528 497
rect 3632 416 3732 497
rect 3880 416 3980 497
rect 3136 403 4084 416
rect 3136 357 3149 403
rect 3571 357 4084 403
rect 3136 344 4084 357
rect 2656 257 2776 301
rect 3136 288 3236 344
rect 150 80 270 124
rect 374 64 494 124
rect 742 112 862 156
rect 966 112 1086 156
rect 1190 64 1310 156
rect 1358 112 1478 156
rect 1670 141 1790 185
rect 1894 152 2014 185
rect 1894 106 1907 152
rect 1953 106 2014 152
rect 2118 141 2238 185
rect 1894 93 2014 106
rect 3116 232 3236 288
rect 3428 232 3548 344
rect 3652 232 3772 344
rect 3964 232 4084 344
rect 374 24 1310 64
rect 2432 24 2552 68
rect 2656 24 2776 68
rect 3116 24 3236 68
rect 3428 24 3548 68
rect 3652 24 3772 68
rect 3964 24 4084 68
<< polycontact >>
rect 1214 632 1260 678
rect 183 366 229 412
rect 387 280 433 326
rect 807 369 853 415
rect 1419 421 1465 467
rect 1218 261 1264 307
rect 1683 300 1729 346
rect 2245 362 2291 408
rect 2493 300 2539 346
rect 2697 421 2743 467
rect 3149 357 3571 403
rect 1907 106 1953 152
<< metal1 >>
rect 0 724 4256 844
rect 95 632 141 645
rect 288 632 356 724
rect 636 647 704 724
rect 288 586 299 632
rect 345 586 356 632
rect 503 632 569 645
rect 141 492 433 518
rect 95 472 433 492
rect 56 412 318 426
rect 56 366 183 412
rect 229 366 318 412
rect 56 354 318 366
rect 387 326 433 472
rect 387 275 433 280
rect 75 229 433 275
rect 549 542 569 632
rect 636 601 647 647
rect 693 601 704 647
rect 766 632 1214 678
rect 1260 632 1271 678
rect 766 542 812 632
rect 1541 586 1609 724
rect 2570 702 2638 724
rect 2570 656 2581 702
rect 2627 656 2638 702
rect 3050 703 3118 724
rect 2700 610 3004 651
rect 2358 609 3004 610
rect 549 496 812 542
rect 884 529 895 575
rect 941 529 1058 575
rect 549 492 569 496
rect 75 204 121 229
rect 503 204 569 492
rect 690 415 878 430
rect 690 369 807 415
rect 853 369 878 415
rect 690 354 878 369
rect 1011 215 1058 529
rect 75 147 121 158
rect 288 137 299 183
rect 345 137 356 183
rect 503 158 523 204
rect 503 147 569 158
rect 656 169 667 215
rect 713 169 724 215
rect 880 169 891 215
rect 937 169 1058 215
rect 1115 513 1126 559
rect 1172 513 1183 559
rect 1541 540 1552 586
rect 1598 540 1609 586
rect 1808 575 1876 586
rect 1115 410 1183 513
rect 1808 529 1818 575
rect 1864 529 1876 575
rect 1808 478 1876 529
rect 1419 467 1876 478
rect 1465 421 1876 467
rect 1419 410 1876 421
rect 1115 364 1356 410
rect 1115 215 1161 364
rect 1310 346 1356 364
rect 1218 307 1264 318
rect 1310 300 1683 346
rect 1729 300 1740 346
rect 1218 254 1264 261
rect 1218 208 1712 254
rect 288 60 356 137
rect 656 60 724 169
rect 1115 158 1161 169
rect 1540 116 1551 162
rect 1597 116 1608 162
rect 1540 60 1608 116
rect 1666 152 1712 208
rect 1808 244 1876 410
rect 1808 198 1819 244
rect 1865 198 1876 244
rect 2032 575 2100 586
rect 2032 529 2043 575
rect 2089 529 2100 575
rect 2358 563 2377 609
rect 2423 605 3004 609
rect 2423 563 2746 605
rect 2032 517 2100 529
rect 2032 471 2754 517
rect 2032 244 2100 471
rect 2686 467 2754 471
rect 2686 421 2697 467
rect 2743 421 2754 467
rect 2818 513 2829 559
rect 2875 513 2886 559
rect 2032 198 2043 244
rect 2089 198 2100 244
rect 2234 362 2245 408
rect 2291 362 2302 408
rect 2234 152 2302 362
rect 2818 403 2886 513
rect 2958 505 3004 605
rect 3050 563 3061 703
rect 3107 563 3118 703
rect 3546 703 3614 724
rect 3165 632 3500 678
rect 3546 657 3557 703
rect 3603 657 3614 703
rect 4102 703 4170 724
rect 3165 505 3211 632
rect 3454 611 3500 632
rect 3660 632 4026 678
rect 3660 611 3706 632
rect 2958 459 3211 505
rect 3298 540 3309 586
rect 3355 540 3368 586
rect 3454 565 3706 611
rect 3298 519 3368 540
rect 3774 540 3785 586
rect 3831 540 3902 586
rect 3774 519 3902 540
rect 3298 449 3902 519
rect 2818 357 3149 403
rect 3571 357 3582 403
rect 2818 346 2898 357
rect 2482 300 2493 346
rect 2539 300 2898 346
rect 3714 311 3902 449
rect 2482 299 2898 300
rect 2830 244 2898 299
rect 1666 106 1907 152
rect 1953 106 2302 152
rect 2349 192 2730 219
rect 2830 198 2841 244
rect 2887 198 2898 244
rect 3298 265 3902 311
rect 3298 244 3366 265
rect 2395 173 2730 192
rect 2349 135 2395 146
rect 2684 152 2730 173
rect 2949 184 3179 230
rect 3298 198 3309 244
rect 3355 198 3366 244
rect 3834 244 3902 265
rect 2949 152 2995 184
rect 2570 81 2581 127
rect 2627 81 2638 127
rect 2684 106 2995 152
rect 3133 152 3179 184
rect 3474 173 3726 219
rect 3834 198 3845 244
rect 3891 198 3902 244
rect 3474 152 3520 173
rect 3041 127 3087 138
rect 2570 60 2638 81
rect 3133 106 3520 152
rect 3680 152 3726 173
rect 3980 152 4026 632
rect 4102 563 4113 703
rect 4159 563 4170 703
rect 3041 60 3087 81
rect 3566 81 3577 127
rect 3623 81 3634 127
rect 3680 106 4026 152
rect 4113 142 4159 153
rect 3566 60 3634 81
rect 4113 60 4159 96
rect 0 -60 4256 60
<< labels >>
flabel metal1 s 690 354 878 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 3774 519 3902 586 0 FreeSans 600 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 724 4256 844 0 FreeSans 600 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 656 183 724 215 0 FreeSans 600 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 56 354 318 426 0 FreeSans 600 0 0 0 CLKN
port 2 nsew clock input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 3298 519 3368 586 1 Q
port 3 nsew default output
rlabel metal1 s 3298 449 3902 519 1 Q
port 3 nsew default output
rlabel metal1 s 3714 311 3902 449 1 Q
port 3 nsew default output
rlabel metal1 s 3298 265 3902 311 1 Q
port 3 nsew default output
rlabel metal1 s 3834 198 3902 265 1 Q
port 3 nsew default output
rlabel metal1 s 3298 198 3366 265 1 Q
port 3 nsew default output
rlabel metal1 s 4102 657 4170 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3546 657 3614 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3050 657 3118 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2570 657 2638 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 657 1609 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 657 704 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 657 356 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4102 656 4170 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3050 656 3118 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2570 656 2638 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 656 1609 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 656 704 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 656 356 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4102 601 4170 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3050 601 3118 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 601 1609 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 601 704 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 601 356 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4102 586 4170 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3050 586 3118 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 586 1609 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 586 356 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4102 563 4170 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3050 563 3118 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 563 1609 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 540 1609 563 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 656 162 724 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 288 162 356 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1540 153 1608 162 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 656 153 724 162 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 288 153 356 162 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 138 4159 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1540 138 1608 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 656 138 724 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 288 138 356 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 127 4159 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3041 127 3087 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1540 127 1608 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 656 127 724 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 288 127 356 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 60 4159 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3566 60 3634 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3041 60 3087 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2570 60 2638 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1540 60 1608 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 656 60 724 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 288 60 356 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string GDS_END 882006
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 873170
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
