magic
tech gf180mcuD
timestamp 1755724134
<< properties >>
string GDS_END 7058056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7057012
<< end >>
