magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< mvnmos >>
rect 124 69 324 333
rect 572 69 772 333
rect 1020 69 1220 333
rect 1468 69 1668 333
rect 1916 69 2116 333
rect 2364 69 2564 333
rect 2812 69 3012 333
rect 3260 69 3460 333
<< mvpmos >>
rect 124 573 324 939
rect 572 573 772 939
rect 1020 573 1220 939
rect 1468 573 1668 939
rect 1916 573 2116 939
rect 2364 573 2564 939
rect 2812 573 3012 939
rect 3260 573 3460 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 324 287 412 333
rect 324 147 353 287
rect 399 147 412 287
rect 324 69 412 147
rect 484 287 572 333
rect 484 147 497 287
rect 543 147 572 287
rect 484 69 572 147
rect 772 287 860 333
rect 772 147 801 287
rect 847 147 860 287
rect 772 69 860 147
rect 932 287 1020 333
rect 932 147 945 287
rect 991 147 1020 287
rect 932 69 1020 147
rect 1220 287 1308 333
rect 1220 147 1249 287
rect 1295 147 1308 287
rect 1220 69 1308 147
rect 1380 287 1468 333
rect 1380 147 1393 287
rect 1439 147 1468 287
rect 1380 69 1468 147
rect 1668 287 1756 333
rect 1668 147 1697 287
rect 1743 147 1756 287
rect 1668 69 1756 147
rect 1828 287 1916 333
rect 1828 147 1841 287
rect 1887 147 1916 287
rect 1828 69 1916 147
rect 2116 287 2204 333
rect 2116 147 2145 287
rect 2191 147 2204 287
rect 2116 69 2204 147
rect 2276 287 2364 333
rect 2276 147 2289 287
rect 2335 147 2364 287
rect 2276 69 2364 147
rect 2564 287 2652 333
rect 2564 147 2593 287
rect 2639 147 2652 287
rect 2564 69 2652 147
rect 2724 287 2812 333
rect 2724 147 2737 287
rect 2783 147 2812 287
rect 2724 69 2812 147
rect 3012 287 3100 333
rect 3012 147 3041 287
rect 3087 147 3100 287
rect 3012 69 3100 147
rect 3172 287 3260 333
rect 3172 147 3185 287
rect 3231 147 3260 287
rect 3172 69 3260 147
rect 3460 287 3548 333
rect 3460 147 3489 287
rect 3535 147 3548 287
rect 3460 69 3548 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 324 861 412 939
rect 324 721 353 861
rect 399 721 412 861
rect 324 573 412 721
rect 484 861 572 939
rect 484 721 497 861
rect 543 721 572 861
rect 484 573 572 721
rect 772 861 860 939
rect 772 721 801 861
rect 847 721 860 861
rect 772 573 860 721
rect 932 861 1020 939
rect 932 721 945 861
rect 991 721 1020 861
rect 932 573 1020 721
rect 1220 861 1308 939
rect 1220 721 1249 861
rect 1295 721 1308 861
rect 1220 573 1308 721
rect 1380 861 1468 939
rect 1380 721 1393 861
rect 1439 721 1468 861
rect 1380 573 1468 721
rect 1668 861 1756 939
rect 1668 721 1697 861
rect 1743 721 1756 861
rect 1668 573 1756 721
rect 1828 861 1916 939
rect 1828 721 1841 861
rect 1887 721 1916 861
rect 1828 573 1916 721
rect 2116 861 2204 939
rect 2116 721 2145 861
rect 2191 721 2204 861
rect 2116 573 2204 721
rect 2276 861 2364 939
rect 2276 721 2289 861
rect 2335 721 2364 861
rect 2276 573 2364 721
rect 2564 861 2652 939
rect 2564 721 2593 861
rect 2639 721 2652 861
rect 2564 573 2652 721
rect 2724 861 2812 939
rect 2724 721 2737 861
rect 2783 721 2812 861
rect 2724 573 2812 721
rect 3012 861 3100 939
rect 3012 721 3041 861
rect 3087 721 3100 861
rect 3012 573 3100 721
rect 3172 861 3260 939
rect 3172 721 3185 861
rect 3231 721 3260 861
rect 3172 573 3260 721
rect 3460 861 3548 939
rect 3460 721 3489 861
rect 3535 721 3548 861
rect 3460 573 3548 721
<< mvndiffc >>
rect 49 147 95 287
rect 353 147 399 287
rect 497 147 543 287
rect 801 147 847 287
rect 945 147 991 287
rect 1249 147 1295 287
rect 1393 147 1439 287
rect 1697 147 1743 287
rect 1841 147 1887 287
rect 2145 147 2191 287
rect 2289 147 2335 287
rect 2593 147 2639 287
rect 2737 147 2783 287
rect 3041 147 3087 287
rect 3185 147 3231 287
rect 3489 147 3535 287
<< mvpdiffc >>
rect 49 721 95 861
rect 353 721 399 861
rect 497 721 543 861
rect 801 721 847 861
rect 945 721 991 861
rect 1249 721 1295 861
rect 1393 721 1439 861
rect 1697 721 1743 861
rect 1841 721 1887 861
rect 2145 721 2191 861
rect 2289 721 2335 861
rect 2593 721 2639 861
rect 2737 721 2783 861
rect 3041 721 3087 861
rect 3185 721 3231 861
rect 3489 721 3535 861
<< polysilicon >>
rect 124 939 324 983
rect 572 939 772 983
rect 1020 939 1220 983
rect 1468 939 1668 983
rect 1916 939 2116 983
rect 2364 939 2564 983
rect 2812 939 3012 983
rect 3260 939 3460 983
rect 124 540 324 573
rect 124 494 265 540
rect 311 494 324 540
rect 124 481 324 494
rect 572 540 772 573
rect 572 494 713 540
rect 759 494 772 540
rect 572 481 772 494
rect 1020 540 1220 573
rect 1020 494 1161 540
rect 1207 494 1220 540
rect 1020 481 1220 494
rect 1468 540 1668 573
rect 1468 494 1609 540
rect 1655 494 1668 540
rect 1468 481 1668 494
rect 1916 540 2116 573
rect 1916 494 2057 540
rect 2103 494 2116 540
rect 1916 481 2116 494
rect 2364 540 2564 573
rect 2364 494 2505 540
rect 2551 494 2564 540
rect 2364 481 2564 494
rect 2812 540 3012 573
rect 2812 494 2953 540
rect 2999 494 3012 540
rect 2812 481 3012 494
rect 3260 540 3460 573
rect 3260 494 3401 540
rect 3447 494 3460 540
rect 3260 481 3460 494
rect 124 412 324 425
rect 124 366 137 412
rect 183 366 324 412
rect 124 333 324 366
rect 572 412 772 425
rect 572 366 585 412
rect 631 366 772 412
rect 572 333 772 366
rect 1020 412 1220 425
rect 1020 366 1033 412
rect 1079 366 1220 412
rect 1020 333 1220 366
rect 1468 412 1668 425
rect 1468 366 1481 412
rect 1527 366 1668 412
rect 1468 333 1668 366
rect 1916 412 2116 425
rect 1916 366 1929 412
rect 1975 366 2116 412
rect 1916 333 2116 366
rect 2364 412 2564 425
rect 2364 366 2377 412
rect 2423 366 2564 412
rect 2364 333 2564 366
rect 2812 412 3012 425
rect 2812 366 2825 412
rect 2871 366 3012 412
rect 2812 333 3012 366
rect 3260 412 3460 425
rect 3260 366 3273 412
rect 3319 366 3460 412
rect 3260 333 3460 366
rect 124 25 324 69
rect 572 25 772 69
rect 1020 25 1220 69
rect 1468 25 1668 69
rect 1916 25 2116 69
rect 2364 25 2564 69
rect 2812 25 3012 69
rect 3260 25 3460 69
<< polycontact >>
rect 265 494 311 540
rect 713 494 759 540
rect 1161 494 1207 540
rect 1609 494 1655 540
rect 2057 494 2103 540
rect 2505 494 2551 540
rect 2953 494 2999 540
rect 3401 494 3447 540
rect 137 366 183 412
rect 585 366 631 412
rect 1033 366 1079 412
rect 1481 366 1527 412
rect 1929 366 1975 412
rect 2377 366 2423 412
rect 2825 366 2871 412
rect 3273 366 3319 412
<< metal1 >>
rect 0 918 3584 1098
rect 49 861 95 872
rect 49 412 95 721
rect 353 861 399 918
rect 353 710 399 721
rect 497 861 543 872
rect 265 540 311 551
rect 49 366 137 412
rect 183 366 194 412
rect 265 298 311 494
rect 497 412 543 721
rect 801 861 847 918
rect 801 710 847 721
rect 945 861 991 872
rect 713 540 759 551
rect 497 366 585 412
rect 631 366 642 412
rect 713 298 759 494
rect 945 412 991 721
rect 1249 861 1295 918
rect 1249 710 1295 721
rect 1393 861 1439 872
rect 1161 540 1207 551
rect 945 366 1033 412
rect 1079 366 1090 412
rect 1161 298 1207 494
rect 1393 412 1439 721
rect 1697 861 1743 918
rect 1697 710 1743 721
rect 1841 861 1887 872
rect 1609 540 1655 551
rect 1393 366 1481 412
rect 1527 366 1538 412
rect 1609 298 1655 494
rect 1841 412 1887 721
rect 2145 861 2191 918
rect 2145 710 2191 721
rect 2289 861 2335 872
rect 2057 540 2103 551
rect 1841 366 1929 412
rect 1975 366 1986 412
rect 2057 298 2103 494
rect 2289 412 2335 721
rect 2593 861 2639 918
rect 2593 710 2639 721
rect 2737 861 2783 872
rect 2505 540 2551 551
rect 2289 366 2377 412
rect 2423 366 2434 412
rect 2505 298 2551 494
rect 2737 412 2783 721
rect 3041 861 3087 918
rect 3041 710 3087 721
rect 3185 861 3231 872
rect 2953 540 2999 551
rect 2737 366 2825 412
rect 2871 366 2882 412
rect 2953 298 2999 494
rect 3185 412 3231 721
rect 3489 861 3535 918
rect 3489 710 3535 721
rect 3401 540 3447 551
rect 3185 366 3273 412
rect 3319 366 3330 412
rect 3401 298 3447 494
rect 49 287 95 298
rect 265 287 399 298
rect 265 252 353 287
rect 49 90 95 147
rect 353 136 399 147
rect 497 287 543 298
rect 713 287 847 298
rect 713 252 801 287
rect 497 90 543 147
rect 801 136 847 147
rect 945 287 991 298
rect 1161 287 1295 298
rect 1161 252 1249 287
rect 945 90 991 147
rect 1249 136 1295 147
rect 1393 287 1439 298
rect 1609 287 1743 298
rect 1609 252 1697 287
rect 1393 90 1439 147
rect 1697 136 1743 147
rect 1841 287 1887 298
rect 2057 287 2191 298
rect 2057 252 2145 287
rect 1841 90 1887 147
rect 2145 136 2191 147
rect 2289 287 2335 298
rect 2505 287 2639 298
rect 2505 252 2593 287
rect 2289 90 2335 147
rect 2593 136 2639 147
rect 2737 287 2783 298
rect 2953 287 3087 298
rect 2953 252 3041 287
rect 2737 90 2783 147
rect 3041 136 3087 147
rect 3185 287 3231 298
rect 3401 287 3535 298
rect 3401 252 3489 287
rect 3185 90 3231 147
rect 3489 136 3535 147
rect 0 -90 3584 90
<< labels >>
flabel metal1 s 0 918 3584 1098 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 3185 90 3231 298 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 3489 710 3535 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3041 710 3087 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2593 710 2639 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2145 710 2191 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 710 1743 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 710 1295 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 710 847 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 710 399 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2737 90 2783 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3584 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string GDS_END 795478
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 785228
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
