magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect 487 1987 1631 2449
rect 263 1986 1631 1987
rect 4 1774 1630 1986
rect 4 1037 1631 1774
rect 4 797 1630 1037
<< mvnmos >>
rect 742 2587 862 2779
rect 1256 2587 1376 2779
rect 518 295 638 659
rect 742 295 862 659
rect 1256 204 1376 658
<< mvpmos >>
rect 742 2116 862 2308
rect 1256 2116 1376 2308
rect 518 939 638 1847
rect 742 939 862 1847
rect 1256 1179 1376 1633
<< mvndiff >>
rect 654 2766 742 2779
rect 654 2720 667 2766
rect 713 2720 742 2766
rect 654 2646 742 2720
rect 654 2600 667 2646
rect 713 2600 742 2646
rect 654 2587 742 2600
rect 862 2766 950 2779
rect 862 2720 891 2766
rect 937 2720 950 2766
rect 862 2646 950 2720
rect 862 2600 891 2646
rect 937 2600 950 2646
rect 862 2587 950 2600
rect 1168 2766 1256 2779
rect 1168 2720 1181 2766
rect 1227 2720 1256 2766
rect 1168 2646 1256 2720
rect 1168 2600 1181 2646
rect 1227 2600 1256 2646
rect 1168 2587 1256 2600
rect 1376 2766 1464 2779
rect 1376 2720 1405 2766
rect 1451 2720 1464 2766
rect 1376 2646 1464 2720
rect 1376 2600 1405 2646
rect 1451 2600 1464 2646
rect 1376 2587 1464 2600
rect 430 646 518 659
rect 430 600 443 646
rect 489 600 518 646
rect 430 500 518 600
rect 430 454 443 500
rect 489 454 518 500
rect 430 354 518 454
rect 430 308 443 354
rect 489 308 518 354
rect 430 295 518 308
rect 638 646 742 659
rect 638 600 667 646
rect 713 600 742 646
rect 638 500 742 600
rect 638 454 667 500
rect 713 454 742 500
rect 638 354 742 454
rect 638 308 667 354
rect 713 308 742 354
rect 638 295 742 308
rect 862 646 950 659
rect 862 600 891 646
rect 937 600 950 646
rect 862 500 950 600
rect 862 454 891 500
rect 937 454 950 500
rect 862 354 950 454
rect 862 308 891 354
rect 937 308 950 354
rect 862 295 950 308
rect 1168 645 1256 658
rect 1168 599 1181 645
rect 1227 599 1256 645
rect 1168 518 1256 599
rect 1168 472 1181 518
rect 1227 472 1256 518
rect 1168 391 1256 472
rect 1168 345 1181 391
rect 1227 345 1256 391
rect 1168 263 1256 345
rect 1168 217 1181 263
rect 1227 217 1256 263
rect 1168 204 1256 217
rect 1376 645 1464 658
rect 1376 599 1405 645
rect 1451 599 1464 645
rect 1376 518 1464 599
rect 1376 472 1405 518
rect 1451 472 1464 518
rect 1376 391 1464 472
rect 1376 345 1405 391
rect 1451 345 1464 391
rect 1376 263 1464 345
rect 1376 217 1405 263
rect 1451 217 1464 263
rect 1376 204 1464 217
<< mvpdiff >>
rect 654 2295 742 2308
rect 654 2249 667 2295
rect 713 2249 742 2295
rect 654 2175 742 2249
rect 654 2129 667 2175
rect 713 2129 742 2175
rect 654 2116 742 2129
rect 862 2295 950 2308
rect 862 2249 891 2295
rect 937 2249 950 2295
rect 862 2175 950 2249
rect 862 2129 891 2175
rect 937 2129 950 2175
rect 862 2116 950 2129
rect 1168 2295 1256 2308
rect 1168 2249 1181 2295
rect 1227 2249 1256 2295
rect 1168 2175 1256 2249
rect 1168 2129 1181 2175
rect 1227 2129 1256 2175
rect 1168 2116 1256 2129
rect 1376 2295 1464 2308
rect 1376 2249 1405 2295
rect 1451 2249 1464 2295
rect 1376 2175 1464 2249
rect 1376 2129 1405 2175
rect 1451 2129 1464 2175
rect 1376 2116 1464 2129
rect 430 1834 518 1847
rect 430 1788 443 1834
rect 489 1788 518 1834
rect 430 1730 518 1788
rect 430 1684 443 1730
rect 489 1684 518 1730
rect 430 1626 518 1684
rect 430 1580 443 1626
rect 489 1580 518 1626
rect 430 1522 518 1580
rect 430 1476 443 1522
rect 489 1476 518 1522
rect 430 1418 518 1476
rect 430 1372 443 1418
rect 489 1372 518 1418
rect 430 1313 518 1372
rect 430 1267 443 1313
rect 489 1267 518 1313
rect 430 1208 518 1267
rect 430 1162 443 1208
rect 489 1162 518 1208
rect 430 1103 518 1162
rect 430 1057 443 1103
rect 489 1057 518 1103
rect 430 998 518 1057
rect 430 952 443 998
rect 489 952 518 998
rect 430 939 518 952
rect 638 1834 742 1847
rect 638 1788 667 1834
rect 713 1788 742 1834
rect 638 1730 742 1788
rect 638 1684 667 1730
rect 713 1684 742 1730
rect 638 1626 742 1684
rect 638 1580 667 1626
rect 713 1580 742 1626
rect 638 1522 742 1580
rect 638 1476 667 1522
rect 713 1476 742 1522
rect 638 1418 742 1476
rect 638 1372 667 1418
rect 713 1372 742 1418
rect 638 1313 742 1372
rect 638 1267 667 1313
rect 713 1267 742 1313
rect 638 1208 742 1267
rect 638 1162 667 1208
rect 713 1162 742 1208
rect 638 1103 742 1162
rect 638 1057 667 1103
rect 713 1057 742 1103
rect 638 998 742 1057
rect 638 952 667 998
rect 713 952 742 998
rect 638 939 742 952
rect 862 1834 950 1847
rect 862 1788 891 1834
rect 937 1788 950 1834
rect 862 1730 950 1788
rect 862 1684 891 1730
rect 937 1684 950 1730
rect 862 1626 950 1684
rect 862 1580 891 1626
rect 937 1580 950 1626
rect 862 1522 950 1580
rect 862 1476 891 1522
rect 937 1476 950 1522
rect 862 1418 950 1476
rect 862 1372 891 1418
rect 937 1372 950 1418
rect 862 1313 950 1372
rect 862 1267 891 1313
rect 937 1267 950 1313
rect 862 1208 950 1267
rect 862 1162 891 1208
rect 937 1162 950 1208
rect 1168 1620 1256 1633
rect 1168 1574 1181 1620
rect 1227 1574 1256 1620
rect 1168 1493 1256 1574
rect 1168 1447 1181 1493
rect 1227 1447 1256 1493
rect 1168 1366 1256 1447
rect 1168 1320 1181 1366
rect 1227 1320 1256 1366
rect 1168 1238 1256 1320
rect 1168 1192 1181 1238
rect 1227 1192 1256 1238
rect 1168 1179 1256 1192
rect 1376 1620 1464 1633
rect 1376 1574 1405 1620
rect 1451 1574 1464 1620
rect 1376 1493 1464 1574
rect 1376 1447 1405 1493
rect 1451 1447 1464 1493
rect 1376 1366 1464 1447
rect 1376 1320 1405 1366
rect 1451 1320 1464 1366
rect 1376 1238 1464 1320
rect 1376 1192 1405 1238
rect 1451 1192 1464 1238
rect 1376 1179 1464 1192
rect 862 1103 950 1162
rect 862 1057 891 1103
rect 937 1057 950 1103
rect 862 998 950 1057
rect 862 952 891 998
rect 937 952 950 998
rect 862 939 950 952
<< mvndiffc >>
rect 667 2720 713 2766
rect 667 2600 713 2646
rect 891 2720 937 2766
rect 891 2600 937 2646
rect 1181 2720 1227 2766
rect 1181 2600 1227 2646
rect 1405 2720 1451 2766
rect 1405 2600 1451 2646
rect 443 600 489 646
rect 443 454 489 500
rect 443 308 489 354
rect 667 600 713 646
rect 667 454 713 500
rect 667 308 713 354
rect 891 600 937 646
rect 891 454 937 500
rect 891 308 937 354
rect 1181 599 1227 645
rect 1181 472 1227 518
rect 1181 345 1227 391
rect 1181 217 1227 263
rect 1405 599 1451 645
rect 1405 472 1451 518
rect 1405 345 1451 391
rect 1405 217 1451 263
<< mvpdiffc >>
rect 667 2249 713 2295
rect 667 2129 713 2175
rect 891 2249 937 2295
rect 891 2129 937 2175
rect 1181 2249 1227 2295
rect 1181 2129 1227 2175
rect 1405 2249 1451 2295
rect 1405 2129 1451 2175
rect 443 1788 489 1834
rect 443 1684 489 1730
rect 443 1580 489 1626
rect 443 1476 489 1522
rect 443 1372 489 1418
rect 443 1267 489 1313
rect 443 1162 489 1208
rect 443 1057 489 1103
rect 443 952 489 998
rect 667 1788 713 1834
rect 667 1684 713 1730
rect 667 1580 713 1626
rect 667 1476 713 1522
rect 667 1372 713 1418
rect 667 1267 713 1313
rect 667 1162 713 1208
rect 667 1057 713 1103
rect 667 952 713 998
rect 891 1788 937 1834
rect 891 1684 937 1730
rect 891 1580 937 1626
rect 891 1476 937 1522
rect 891 1372 937 1418
rect 891 1267 937 1313
rect 891 1162 937 1208
rect 1181 1574 1227 1620
rect 1181 1447 1227 1493
rect 1181 1320 1227 1366
rect 1181 1192 1227 1238
rect 1405 1574 1451 1620
rect 1405 1447 1451 1493
rect 1405 1320 1451 1366
rect 1405 1192 1451 1238
rect 891 1057 937 1103
rect 891 952 937 998
<< psubdiff >>
rect 149 2775 466 2834
rect 149 2729 205 2775
rect 251 2729 363 2775
rect 409 2729 466 2775
rect 149 2669 466 2729
rect 110 508 243 567
rect 110 462 153 508
rect 199 462 243 508
rect 110 345 243 462
rect 110 299 153 345
rect 199 299 243 345
rect 110 239 243 299
<< nsubdiff >>
rect 110 1801 243 1846
rect 110 1755 153 1801
rect 199 1755 243 1801
rect 110 1608 243 1755
rect 110 1562 153 1608
rect 199 1562 243 1608
rect 110 1415 243 1562
rect 110 1369 153 1415
rect 199 1369 243 1415
rect 110 1223 243 1369
rect 110 1177 153 1223
rect 199 1177 243 1223
rect 110 1015 243 1177
<< psubdiffcont >>
rect 205 2729 251 2775
rect 363 2729 409 2775
rect 153 462 199 508
rect 153 299 199 345
<< nsubdiffcont >>
rect 153 1755 199 1801
rect 153 1562 199 1608
rect 153 1369 199 1415
rect 153 1177 199 1223
<< polysilicon >>
rect 742 2779 862 2823
rect 1256 2779 1376 2823
rect 742 2308 862 2587
rect 1256 2527 1376 2587
rect 1582 2527 1666 2528
rect 1256 2509 1666 2527
rect 1256 2461 1601 2509
rect 1257 2352 1375 2381
rect 1582 2369 1601 2461
rect 1647 2369 1666 2509
rect 1256 2308 1376 2352
rect 375 2091 459 2110
rect 375 2045 394 2091
rect 440 2056 459 2091
rect 742 2056 862 2116
rect 440 2045 862 2056
rect 375 1996 862 2045
rect 1256 2028 1376 2116
rect 1256 2009 1439 2028
rect 1256 1963 1374 2009
rect 1420 1963 1439 2009
rect 1256 1944 1439 1963
rect 519 1891 637 1918
rect 743 1891 861 1918
rect 518 1847 638 1891
rect 742 1847 862 1891
rect 1582 1762 1666 2369
rect 1256 1693 1666 1762
rect 1256 1633 1376 1693
rect 1256 1135 1376 1179
rect 1256 1105 1375 1135
rect 518 864 638 939
rect 742 864 862 939
rect 518 819 1024 864
rect 518 773 904 819
rect 950 773 1024 819
rect 1490 835 1683 880
rect 1490 804 1563 835
rect 1489 803 1563 804
rect 518 727 1024 773
rect 1256 789 1563 803
rect 1609 789 1683 835
rect 1256 743 1683 789
rect 518 659 638 727
rect 742 659 862 727
rect 1256 658 1376 743
rect 518 251 638 295
rect 742 251 862 295
rect 519 221 637 251
rect 743 221 861 251
rect 1256 160 1376 204
rect 1256 130 1375 160
<< polycontact >>
rect 1601 2369 1647 2509
rect 394 2045 440 2091
rect 1374 1963 1420 2009
rect 904 773 950 819
rect 1563 789 1609 835
<< metal1 >>
rect 632 2864 1472 2968
rect 158 2775 457 2825
rect 158 2771 205 2775
rect 113 2731 205 2771
rect 113 2679 150 2731
rect 202 2729 205 2731
rect 251 2729 363 2775
rect 409 2729 457 2775
rect 202 2679 457 2729
rect 113 2678 457 2679
rect 632 2766 748 2864
rect 891 2771 937 2779
rect 632 2720 667 2766
rect 713 2720 748 2766
rect 113 2513 240 2678
rect 113 2461 150 2513
rect 202 2461 240 2513
rect 113 2420 240 2461
rect 632 2646 748 2720
rect 632 2600 667 2646
rect 713 2600 748 2646
rect 632 2295 748 2600
rect 851 2766 978 2771
rect 851 2731 891 2766
rect 937 2731 978 2766
rect 851 2679 888 2731
rect 940 2679 978 2731
rect 851 2646 978 2679
rect 851 2600 891 2646
rect 937 2600 978 2646
rect 1181 2766 1227 2779
rect 1181 2646 1227 2720
rect 851 2513 978 2600
rect 851 2461 888 2513
rect 940 2461 978 2513
rect 851 2420 978 2461
rect 1146 2600 1181 2628
rect 1370 2766 1472 2864
rect 1370 2720 1405 2766
rect 1451 2720 1472 2766
rect 1370 2646 1472 2720
rect 1227 2600 1262 2628
rect 632 2249 667 2295
rect 713 2249 748 2295
rect 632 2175 748 2249
rect 632 2129 667 2175
rect 713 2129 748 2175
rect 632 2116 748 2129
rect 856 2295 972 2308
rect 856 2249 891 2295
rect 937 2249 972 2295
rect 856 2175 972 2249
rect 856 2129 891 2175
rect 937 2129 972 2175
rect 383 2091 451 2102
rect 383 2045 394 2091
rect 440 2045 451 2091
rect 383 2039 451 2045
rect 359 2038 480 2039
rect 359 1946 748 2038
rect 443 1837 489 1847
rect 119 1834 524 1837
rect 119 1801 443 1834
rect 119 1755 153 1801
rect 199 1788 443 1801
rect 489 1788 524 1834
rect 199 1772 524 1788
rect 119 1720 156 1755
rect 208 1730 524 1772
rect 208 1720 443 1730
rect 119 1684 443 1720
rect 489 1684 524 1730
rect 119 1626 524 1684
rect 119 1608 443 1626
rect 119 1562 153 1608
rect 199 1580 443 1608
rect 489 1580 524 1626
rect 199 1562 524 1580
rect 119 1554 524 1562
rect 119 1502 156 1554
rect 208 1522 524 1554
rect 208 1502 443 1522
rect 119 1476 443 1502
rect 489 1476 524 1522
rect 119 1418 524 1476
rect 119 1415 443 1418
rect 119 1369 153 1415
rect 199 1372 443 1415
rect 489 1372 524 1418
rect 199 1369 524 1372
rect 119 1336 524 1369
rect 119 1284 156 1336
rect 208 1313 524 1336
rect 208 1284 443 1313
rect 119 1267 443 1284
rect 489 1267 524 1313
rect 119 1223 524 1267
rect 119 1177 153 1223
rect 199 1208 524 1223
rect 199 1177 443 1208
rect 119 1162 443 1177
rect 489 1162 524 1208
rect 119 1103 524 1162
rect 119 1057 443 1103
rect 489 1057 524 1103
rect 119 998 524 1057
rect 119 952 443 998
rect 489 952 524 998
rect 119 947 524 952
rect 632 1834 748 1946
rect 856 1916 972 2129
rect 1146 2295 1262 2600
rect 1146 2249 1181 2295
rect 1227 2249 1262 2295
rect 1146 2175 1262 2249
rect 1146 2129 1181 2175
rect 1227 2129 1262 2175
rect 632 1788 667 1834
rect 713 1788 748 1834
rect 632 1730 748 1788
rect 632 1684 667 1730
rect 713 1684 748 1730
rect 632 1626 748 1684
rect 632 1580 667 1626
rect 713 1580 748 1626
rect 632 1522 748 1580
rect 632 1476 667 1522
rect 713 1476 748 1522
rect 632 1418 748 1476
rect 632 1372 667 1418
rect 713 1372 748 1418
rect 632 1313 748 1372
rect 632 1267 667 1313
rect 713 1267 748 1313
rect 632 1208 748 1267
rect 632 1162 667 1208
rect 713 1162 748 1208
rect 632 1103 748 1162
rect 850 1876 978 1916
rect 850 1824 888 1876
rect 940 1824 978 1876
rect 850 1788 891 1824
rect 937 1788 978 1824
rect 850 1730 978 1788
rect 850 1684 891 1730
rect 937 1684 978 1730
rect 850 1658 978 1684
rect 850 1606 888 1658
rect 940 1606 978 1658
rect 850 1580 891 1606
rect 937 1580 978 1606
rect 850 1522 978 1580
rect 850 1476 891 1522
rect 937 1476 978 1522
rect 850 1440 978 1476
rect 850 1388 888 1440
rect 940 1388 978 1440
rect 850 1372 891 1388
rect 937 1372 978 1388
rect 850 1313 978 1372
rect 850 1267 891 1313
rect 937 1267 978 1313
rect 850 1222 978 1267
rect 850 1170 888 1222
rect 940 1170 978 1222
rect 850 1162 891 1170
rect 937 1162 978 1170
rect 850 1130 978 1162
rect 1146 1620 1262 2129
rect 1370 2600 1405 2646
rect 1451 2600 1472 2646
rect 1370 2295 1472 2600
rect 1370 2249 1405 2295
rect 1451 2249 1472 2295
rect 1370 2175 1472 2249
rect 1565 2558 1692 2598
rect 1565 2509 1602 2558
rect 1565 2369 1601 2509
rect 1654 2506 1692 2558
rect 1647 2369 1692 2506
rect 1565 2340 1692 2369
rect 1565 2288 1602 2340
rect 1654 2288 1692 2340
rect 1565 2247 1692 2288
rect 1370 2129 1405 2175
rect 1451 2129 1472 2175
rect 1370 2116 1472 2129
rect 1340 2009 1691 2045
rect 1340 1963 1374 2009
rect 1420 2005 1691 2009
rect 1420 1963 1601 2005
rect 1340 1953 1601 1963
rect 1653 1953 1691 2005
rect 1340 1926 1691 1953
rect 1564 1787 1691 1926
rect 1564 1735 1601 1787
rect 1653 1735 1691 1787
rect 1564 1694 1691 1735
rect 1146 1574 1181 1620
rect 1227 1574 1262 1620
rect 1146 1493 1262 1574
rect 1146 1447 1181 1493
rect 1227 1447 1262 1493
rect 1146 1366 1262 1447
rect 1146 1320 1181 1366
rect 1227 1320 1262 1366
rect 1146 1238 1262 1320
rect 1146 1192 1181 1238
rect 1227 1192 1262 1238
rect 632 1057 667 1103
rect 713 1057 748 1103
rect 632 998 748 1057
rect 632 952 667 998
rect 713 952 748 998
rect 443 939 489 947
rect 443 649 489 659
rect 115 646 524 649
rect 115 609 443 646
rect 115 557 152 609
rect 204 600 443 609
rect 489 600 524 646
rect 204 557 524 600
rect 115 508 524 557
rect 632 646 748 952
rect 891 1103 937 1130
rect 891 998 937 1057
rect 891 939 937 952
rect 1146 855 1262 1192
rect 870 819 1262 855
rect 870 773 904 819
rect 950 773 1262 819
rect 870 736 1262 773
rect 1145 735 1262 736
rect 891 649 937 659
rect 632 600 667 646
rect 713 600 748 646
rect 632 539 748 600
rect 851 646 978 649
rect 851 609 891 646
rect 937 609 978 646
rect 851 557 888 609
rect 940 557 978 609
rect 1146 645 1262 735
rect 1146 599 1181 645
rect 1227 599 1262 645
rect 1146 561 1262 599
rect 1340 1620 1451 1633
rect 1340 1574 1405 1620
rect 1340 1493 1451 1574
rect 1340 1447 1405 1493
rect 1340 1366 1451 1447
rect 1340 1320 1405 1366
rect 1340 1238 1451 1320
rect 1340 1192 1405 1238
rect 1340 1179 1451 1192
rect 1340 658 1450 1179
rect 1564 871 1644 1694
rect 1529 835 1644 871
rect 1529 789 1563 835
rect 1609 789 1644 835
rect 1529 752 1644 789
rect 1340 645 1451 658
rect 1340 599 1405 645
rect 1340 563 1451 599
rect 115 462 153 508
rect 199 500 524 508
rect 199 462 443 500
rect 115 454 443 462
rect 489 454 524 500
rect 667 500 713 539
rect 115 391 524 454
rect 115 339 152 391
rect 204 354 524 391
rect 204 339 443 354
rect 115 299 153 339
rect 199 308 443 339
rect 489 308 524 354
rect 632 454 667 473
rect 851 500 978 557
rect 713 454 748 473
rect 632 354 748 454
rect 632 353 667 354
rect 199 303 524 308
rect 713 353 748 354
rect 851 454 891 500
rect 937 454 978 500
rect 851 391 978 454
rect 199 299 242 303
rect 115 298 242 299
rect 119 248 234 298
rect 443 295 489 303
rect 667 295 713 308
rect 851 339 888 391
rect 940 339 978 391
rect 851 308 891 339
rect 937 308 978 339
rect 851 298 978 308
rect 1181 518 1227 561
rect 1181 391 1227 472
rect 891 295 937 298
rect 1181 263 1227 345
rect 1181 204 1227 217
rect 1340 523 1485 563
rect 1340 471 1395 523
rect 1447 518 1485 523
rect 1451 472 1485 518
rect 1447 471 1485 472
rect 1340 391 1485 471
rect 1340 345 1405 391
rect 1451 345 1485 391
rect 1340 305 1485 345
rect 1340 253 1395 305
rect 1447 263 1485 305
rect 1340 217 1405 253
rect 1451 217 1485 263
rect 1340 212 1485 217
rect 1405 204 1451 212
<< via1 >>
rect 150 2679 202 2731
rect 150 2461 202 2513
rect 888 2720 891 2731
rect 891 2720 937 2731
rect 937 2720 940 2731
rect 888 2679 940 2720
rect 888 2461 940 2513
rect 156 1755 199 1772
rect 199 1755 208 1772
rect 156 1720 208 1755
rect 156 1502 208 1554
rect 156 1284 208 1336
rect 888 1834 940 1876
rect 888 1824 891 1834
rect 891 1824 937 1834
rect 937 1824 940 1834
rect 888 1626 940 1658
rect 888 1606 891 1626
rect 891 1606 937 1626
rect 937 1606 940 1626
rect 888 1418 940 1440
rect 888 1388 891 1418
rect 891 1388 937 1418
rect 937 1388 940 1418
rect 888 1208 940 1222
rect 888 1170 891 1208
rect 891 1170 937 1208
rect 937 1170 940 1208
rect 1602 2509 1654 2558
rect 1602 2506 1647 2509
rect 1647 2506 1654 2509
rect 1602 2288 1654 2340
rect 1601 1953 1653 2005
rect 1601 1735 1653 1787
rect 152 557 204 609
rect 888 600 891 609
rect 891 600 937 609
rect 937 600 940 609
rect 888 557 940 600
rect 152 345 204 391
rect 152 339 153 345
rect 153 339 199 345
rect 199 339 204 345
rect 888 354 940 391
rect 888 339 891 354
rect 891 339 937 354
rect 937 339 940 354
rect 1395 518 1447 523
rect 1395 472 1405 518
rect 1405 472 1447 518
rect 1395 471 1447 472
rect 1395 263 1447 305
rect 1395 253 1405 263
rect 1405 253 1447 263
<< metal2 >>
rect 113 2842 240 2880
rect 113 2786 148 2842
rect 204 2786 240 2842
rect 113 2731 240 2786
rect 113 2679 150 2731
rect 202 2679 240 2731
rect 113 2624 240 2679
rect 113 2568 148 2624
rect 204 2568 240 2624
rect 113 2513 240 2568
rect 113 2461 150 2513
rect 202 2461 240 2513
rect 113 2406 240 2461
rect 113 2350 148 2406
rect 204 2350 240 2406
rect 113 2312 240 2350
rect 851 2842 978 2880
rect 851 2786 886 2842
rect 942 2786 978 2842
rect 851 2731 978 2786
rect 851 2679 888 2731
rect 940 2679 978 2731
rect 851 2624 978 2679
rect 851 2568 886 2624
rect 942 2568 978 2624
rect 851 2513 978 2568
rect 851 2461 888 2513
rect 940 2461 978 2513
rect 851 2406 978 2461
rect 851 2350 886 2406
rect 942 2350 978 2406
rect 851 2312 978 2350
rect 1565 2558 1692 2598
rect 1565 2506 1602 2558
rect 1654 2506 1692 2558
rect 1565 2340 1692 2506
rect 1565 2288 1602 2340
rect 1654 2288 1692 2340
rect 1565 2247 1692 2288
rect 1564 2005 1691 2045
rect 1564 1953 1601 2005
rect 1653 1953 1691 2005
rect 850 1878 978 1916
rect 850 1822 886 1878
rect 942 1822 978 1878
rect 119 1774 247 1812
rect 119 1718 154 1774
rect 210 1718 247 1774
rect 119 1556 247 1718
rect 119 1500 154 1556
rect 210 1500 247 1556
rect 119 1338 247 1500
rect 119 1282 154 1338
rect 210 1282 247 1338
rect 119 1244 247 1282
rect 850 1660 978 1822
rect 1564 1787 1691 1953
rect 1564 1735 1601 1787
rect 1653 1735 1691 1787
rect 1564 1694 1691 1735
rect 850 1604 886 1660
rect 942 1604 978 1660
rect 850 1442 978 1604
rect 850 1386 886 1442
rect 942 1386 978 1442
rect 850 1224 978 1386
rect 850 1168 886 1224
rect 942 1168 978 1224
rect 850 1130 978 1168
rect 114 611 242 649
rect 114 555 150 611
rect 206 555 242 611
rect 114 393 242 555
rect 114 337 150 393
rect 206 337 242 393
rect 114 298 242 337
rect 850 611 978 649
rect 850 555 886 611
rect 942 555 978 611
rect 850 393 978 555
rect 850 337 886 393
rect 942 337 978 393
rect 850 298 978 337
rect 1358 523 1485 563
rect 1358 471 1395 523
rect 1447 471 1485 523
rect 1358 305 1485 471
rect 1358 253 1395 305
rect 1447 253 1485 305
rect 1358 212 1485 253
<< via2 >>
rect 148 2786 204 2842
rect 148 2568 204 2624
rect 148 2350 204 2406
rect 886 2786 942 2842
rect 886 2568 942 2624
rect 886 2350 942 2406
rect 886 1876 942 1878
rect 886 1824 888 1876
rect 888 1824 940 1876
rect 940 1824 942 1876
rect 886 1822 942 1824
rect 154 1772 210 1774
rect 154 1720 156 1772
rect 156 1720 208 1772
rect 208 1720 210 1772
rect 154 1718 210 1720
rect 154 1554 210 1556
rect 154 1502 156 1554
rect 156 1502 208 1554
rect 208 1502 210 1554
rect 154 1500 210 1502
rect 154 1336 210 1338
rect 154 1284 156 1336
rect 156 1284 208 1336
rect 208 1284 210 1336
rect 154 1282 210 1284
rect 886 1658 942 1660
rect 886 1606 888 1658
rect 888 1606 940 1658
rect 940 1606 942 1658
rect 886 1604 942 1606
rect 886 1440 942 1442
rect 886 1388 888 1440
rect 888 1388 940 1440
rect 940 1388 942 1440
rect 886 1386 942 1388
rect 886 1222 942 1224
rect 886 1170 888 1222
rect 888 1170 940 1222
rect 940 1170 942 1222
rect 886 1168 942 1170
rect 150 609 206 611
rect 150 557 152 609
rect 152 557 204 609
rect 204 557 206 609
rect 150 555 206 557
rect 150 391 206 393
rect 150 339 152 391
rect 152 339 204 391
rect 204 339 206 391
rect 150 337 206 339
rect 886 609 942 611
rect 886 557 888 609
rect 888 557 940 609
rect 940 557 942 609
rect 886 555 942 557
rect 886 391 942 393
rect 886 339 888 391
rect 888 339 940 391
rect 940 339 942 391
rect 886 337 942 339
<< metal3 >>
rect -1 2842 1692 2916
rect -1 2786 148 2842
rect 204 2786 886 2842
rect 942 2786 1692 2842
rect -1 2624 1692 2786
rect -1 2568 148 2624
rect 204 2568 886 2624
rect 942 2568 1692 2624
rect -1 2406 1692 2568
rect -1 2350 148 2406
rect 204 2350 886 2406
rect 942 2350 1692 2406
rect -1 2234 1692 2350
rect -1 1878 1692 1986
rect -1 1822 886 1878
rect 942 1822 1692 1878
rect -1 1774 1692 1822
rect -1 1718 154 1774
rect 210 1718 1692 1774
rect -1 1660 1692 1718
rect -1 1604 886 1660
rect 942 1604 1692 1660
rect -1 1556 1692 1604
rect -1 1500 154 1556
rect 210 1500 1692 1556
rect -1 1442 1692 1500
rect -1 1386 886 1442
rect 942 1386 1692 1442
rect -1 1338 1692 1386
rect -1 1282 154 1338
rect 210 1282 1692 1338
rect -1 1224 1692 1282
rect -1 1168 886 1224
rect 942 1168 1692 1224
rect -1 1078 1692 1168
rect -90 611 1692 907
rect -90 555 150 611
rect 206 555 886 611
rect 942 555 1692 611
rect -90 393 1692 555
rect -90 337 150 393
rect 206 337 886 393
rect 942 337 1692 393
rect -90 -1 1692 337
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_0
timestamp 1755724134
transform 1 0 927 0 1 796
box 0 0 1 1
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_1
timestamp 1755724134
transform 1 0 1586 0 1 812
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1755724134
transform 1 0 1624 0 1 2439
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1755724134
transform 1 0 1397 0 1 1986
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1755724134
transform 1 0 417 0 1 2068
box 0 0 1 1
use M1_PSUB$$45110316_512x8m81  M1_PSUB$$45110316_512x8m81_0
timestamp 1755724134
transform 1 0 307 0 1 2752
box 0 0 1 1
use M2_M1$$43379756_153_512x8m81  M2_M1$$43379756_153_512x8m81_0
timestamp 1755724134
transform 1 0 914 0 1 1523
box 0 0 1 1
use M2_M1$$43380780_152_512x8m81  M2_M1$$43380780_152_512x8m81_0
timestamp 1755724134
transform 1 0 182 0 1 1528
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_0
timestamp 1755724134
transform 1 0 1628 0 1 2423
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_1
timestamp 1755724134
transform 1 0 1627 0 1 1870
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_2
timestamp 1755724134
transform 1 0 1421 0 1 388
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_3
timestamp 1755724134
transform 1 0 178 0 1 474
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_4
timestamp 1755724134
transform 1 0 914 0 1 2596
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_5
timestamp 1755724134
transform 1 0 176 0 1 2596
box 0 0 1 1
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_6
timestamp 1755724134
transform 1 0 914 0 1 474
box 0 0 1 1
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_0
timestamp 1755724134
transform 1 0 914 0 1 474
box 0 0 1 1
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_1
timestamp 1755724134
transform 1 0 178 0 1 474
box 0 0 1 1
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_0
timestamp 1755724134
transform 1 0 182 0 1 1528
box 0 0 1 1
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_1
timestamp 1755724134
transform 1 0 176 0 1 2596
box 0 0 1 1
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_2
timestamp 1755724134
transform 1 0 914 0 1 2596
box 0 0 1 1
use M3_M2$$47333420_150_512x8m81  M3_M2$$47333420_150_512x8m81_0
timestamp 1755724134
transform 1 0 914 0 1 1523
box 0 0 1 1
use nmos_1p2$$47329324_512x8m81  nmos_1p2$$47329324_512x8m81_0
timestamp 1755724134
transform 1 0 549 0 1 295
box -31 0 -30 1
use nmos_1p2_157_512x8m81  nmos_1p2_157_512x8m81_0
timestamp 1755724134
transform 1 0 1287 0 1 204
box -31 0 -30 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1755724134
transform 1 0 742 0 -1 2779
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1755724134
transform 1 0 1256 0 -1 2779
box 0 0 1 1
use pmos_1p2$$47331372_512x8m81  pmos_1p2$$47331372_512x8m81_0
timestamp 1755724134
transform 1 0 549 0 1 939
box -31 0 -30 1
use pmos_1p2_160_512x8m81  pmos_1p2_160_512x8m81_0
timestamp 1755724134
transform 1 0 1287 0 1 1179
box -31 0 -30 1
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_0
timestamp 1755724134
transform 1 0 1287 0 -1 2308
box -31 0 -30 1
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_1
timestamp 1755724134
transform 1 0 773 0 -1 2308
box -31 0 -30 1
<< labels >>
rlabel metal3 s 202 2584 202 2584 4 vss
port 1 nsew
rlabel metal3 s 132 367 132 367 4 vss
port 1 nsew
rlabel metal3 s 156 1498 156 1498 4 vdd
port 2 nsew
rlabel metal1 s 1627 2462 1627 2462 4 enb
port 3 nsew
rlabel metal1 s 1632 1789 1632 1789 4 en
port 4 nsew
rlabel metal1 s 690 413 690 413 4 ab
port 5 nsew
rlabel metal1 s 1416 413 1416 413 4 a
port 6 nsew
<< properties >>
string GDS_END 203968
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 199664
<< end >>
