magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< polysilicon >>
rect 803 8977 1033 8996
rect 803 8931 845 8977
rect 985 8931 1033 8977
rect 803 8900 1033 8931
rect 2677 8977 2907 8996
rect 2677 8931 2719 8977
rect 2859 8931 2907 8977
rect 2677 8900 2907 8931
rect 3151 8977 3381 8996
rect 3151 8931 3193 8977
rect 3333 8931 3381 8977
rect 3151 8900 3381 8931
rect 5025 8977 5255 8996
rect 5025 8931 5067 8977
rect 5207 8931 5255 8977
rect 5025 8900 5255 8931
rect 5499 8977 5729 8996
rect 5499 8931 5541 8977
rect 5681 8931 5729 8977
rect 5499 8900 5729 8931
rect 7373 8977 7603 8996
rect 7373 8931 7415 8977
rect 7555 8931 7603 8977
rect 7373 8900 7603 8931
rect 7847 8977 8077 8996
rect 7847 8931 7894 8977
rect 8034 8931 8077 8977
rect 7847 8900 8077 8931
rect 9721 8977 9951 8996
rect 9721 8931 9767 8977
rect 9907 8931 9951 8977
rect 9721 8900 9951 8931
rect 803 1105 1033 1124
rect 803 1059 845 1105
rect 985 1059 1033 1105
rect 803 1028 1033 1059
rect 2677 1105 2907 1124
rect 2677 1059 2719 1105
rect 2859 1059 2907 1105
rect 2677 1028 2907 1059
rect 3151 1105 3381 1124
rect 3151 1059 3193 1105
rect 3333 1059 3381 1105
rect 3151 1028 3381 1059
rect 5025 1105 5255 1124
rect 5025 1059 5067 1105
rect 5207 1059 5255 1105
rect 5025 1028 5255 1059
rect 5499 1105 5729 1124
rect 5499 1059 5541 1105
rect 5681 1059 5729 1105
rect 5499 1028 5729 1059
rect 7373 1105 7603 1124
rect 7373 1059 7415 1105
rect 7555 1059 7603 1105
rect 7373 1028 7603 1059
rect 7847 1105 8077 1124
rect 7847 1059 7894 1105
rect 8034 1059 8077 1105
rect 7847 1028 8077 1059
rect 9721 1105 9951 1124
rect 9721 1059 9767 1105
rect 9907 1059 9951 1105
rect 9721 1028 9951 1059
<< polycontact >>
rect 845 8931 985 8977
rect 2719 8931 2859 8977
rect 3193 8931 3333 8977
rect 5067 8931 5207 8977
rect 5541 8931 5681 8977
rect 7415 8931 7555 8977
rect 7894 8931 8034 8977
rect 9767 8931 9907 8977
rect 845 1059 985 1105
rect 2719 1059 2859 1105
rect 3193 1059 3333 1105
rect 5067 1059 5207 1105
rect 5541 1059 5681 1105
rect 7415 1059 7555 1105
rect 7894 1059 8034 1105
rect 9767 1059 9907 1105
<< metal1 >>
rect -440 9400 5218 9508
rect -440 9240 3344 9340
rect -440 9080 2870 9180
rect -440 8977 996 9020
rect -440 8931 845 8977
rect 985 8931 996 8977
rect -440 8920 996 8931
rect 2708 8977 2870 9080
rect 2708 8931 2719 8977
rect 2859 8931 2870 8977
rect 2708 8920 2870 8931
rect 3182 8977 3344 9240
rect 3182 8931 3193 8977
rect 3333 8931 3344 8977
rect 3182 8920 3344 8931
rect 5056 8977 5218 9400
rect 5532 9400 11180 9508
rect 5532 8988 5694 9400
rect 7404 9240 11180 9340
rect 5056 8931 5067 8977
rect 5207 8931 5218 8977
rect 5056 8920 5218 8931
rect 5530 8977 5692 8988
rect 5530 8931 5541 8977
rect 5681 8931 5692 8977
rect 5530 8920 5692 8931
rect 7404 8977 7566 9240
rect 7404 8931 7415 8977
rect 7555 8931 7566 8977
rect 7404 8920 7566 8931
rect 7883 9080 11180 9180
rect 7883 8977 8045 9080
rect 7883 8931 7894 8977
rect 8034 8931 8045 8977
rect 7883 8920 8045 8931
rect 9756 8977 11180 9020
rect 9756 8931 9767 8977
rect 9907 8931 11180 8977
rect 9756 8920 11180 8931
rect 893 1116 939 8920
rect 2772 1116 2818 8920
rect 3242 1116 3288 8920
rect 5114 1116 5160 8920
rect 5588 1116 5634 8920
rect 7462 1116 7508 8920
rect 7941 1116 7987 8920
rect 9814 1116 9860 8920
rect 834 1105 996 1116
rect 834 1059 845 1105
rect 985 1059 996 1105
rect 834 1048 996 1059
rect 2708 1105 2870 1116
rect 2708 1059 2719 1105
rect 2859 1059 2870 1105
rect 2708 1048 2870 1059
rect 3182 1105 3344 1116
rect 3182 1059 3193 1105
rect 3333 1059 3344 1105
rect 3182 1048 3344 1059
rect 5056 1105 5218 1116
rect 5056 1059 5067 1105
rect 5207 1059 5218 1105
rect 5056 1048 5218 1059
rect 5530 1105 5692 1116
rect 5530 1059 5541 1105
rect 5681 1059 5692 1105
rect 5530 1048 5692 1059
rect 7404 1105 7566 1116
rect 7404 1059 7415 1105
rect 7555 1059 7566 1105
rect 7404 1048 7566 1059
rect 7883 1105 8045 1116
rect 7883 1059 7894 1105
rect 8034 1059 8045 1105
rect 7883 1048 8045 1059
rect 9756 1105 9918 1116
rect 9756 1059 9767 1105
rect 9907 1059 9918 1105
rect 9756 1048 9918 1059
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_0
timestamp 1755724134
transform 1 0 7641 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_1
timestamp 1755724134
transform 1 0 5293 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_2
timestamp 1755724134
transform 1 0 2945 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_3
timestamp 1755724134
transform 1 0 597 0 1 680
box 48 444 2468 8220
use GR_NMOS_4T  GR_NMOS_4T_0
timestamp 1755724134
transform 1 0 363 0 1 436
box -1730 -583 11766 10481
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1755724134
transform 0 1 5137 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1755724134
transform 0 1 5137 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1755724134
transform 0 1 915 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_3
timestamp 1755724134
transform 0 1 3263 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_4
timestamp 1755724134
transform 0 1 9837 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_5
timestamp 1755724134
transform 0 1 915 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_6
timestamp 1755724134
transform 0 1 7964 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_7
timestamp 1755724134
transform 0 1 5611 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_8
timestamp 1755724134
transform 0 1 7485 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_9
timestamp 1755724134
transform 0 1 2789 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_10
timestamp 1755724134
transform 0 1 3263 1 0 8954
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_11
timestamp 1755724134
transform 0 1 5611 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_12
timestamp 1755724134
transform 0 1 7485 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_13
timestamp 1755724134
transform 0 1 7964 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_14
timestamp 1755724134
transform 0 1 9837 1 0 1082
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_15
timestamp 1755724134
transform 0 1 2789 1 0 1082
box 0 0 1 1
use nmos_4T_metal_stack  nmos_4T_metal_stack_0
timestamp 1755724134
transform -1 0 10151 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_1
timestamp 1755724134
transform 1 0 2951 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_2
timestamp 1755724134
transform 1 0 5299 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_3
timestamp 1755724134
transform 1 0 7647 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_4
timestamp 1755724134
transform 1 0 603 0 1 812
box -44 400 2074 8000
<< properties >>
string GDS_END 3548710
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3542578
string path 199.100 223.150 199.100 26.975 
<< end >>
