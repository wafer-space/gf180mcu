magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< psubdiff >>
rect 0 69946 1000 69968
rect 0 69897 178 69946
rect 0 13151 25 69897
rect 71 69800 178 69897
rect 824 69897 1000 69946
rect 824 69800 929 69897
rect 71 69778 929 69800
rect 71 13287 93 69778
rect 907 13287 929 69778
rect 71 13265 929 13287
rect 71 13151 178 13265
rect 0 13119 178 13151
rect 824 13151 929 13265
rect 975 13151 1000 69897
rect 824 13119 1000 13151
rect 0 13097 1000 13119
<< psubdiffcont >>
rect 25 13151 71 69897
rect 178 69800 824 69946
rect 178 13119 824 13265
rect 929 13151 975 69897
<< metal1 >>
rect -32 69946 1032 69957
rect -32 69897 178 69946
rect -32 13151 25 69897
rect 71 69800 178 69897
rect 824 69897 1032 69946
rect 824 69800 929 69897
rect 71 69789 929 69800
rect 71 64954 82 69789
rect 918 64954 929 69789
rect 71 64822 929 64954
rect 71 64770 232 64822
rect 284 64770 356 64822
rect 408 64770 480 64822
rect 532 64770 604 64822
rect 656 64770 728 64822
rect 780 64770 929 64822
rect 71 64698 929 64770
rect 71 64646 232 64698
rect 284 64646 356 64698
rect 408 64646 480 64698
rect 532 64646 604 64698
rect 656 64646 728 64698
rect 780 64646 929 64698
rect 71 64574 929 64646
rect 71 64522 232 64574
rect 284 64522 356 64574
rect 408 64522 480 64574
rect 532 64522 604 64574
rect 656 64522 728 64574
rect 780 64522 929 64574
rect 71 64450 929 64522
rect 71 64398 232 64450
rect 284 64398 356 64450
rect 408 64398 480 64450
rect 532 64398 604 64450
rect 656 64398 728 64450
rect 780 64398 929 64450
rect 71 64326 929 64398
rect 71 64274 232 64326
rect 284 64274 356 64326
rect 408 64274 480 64326
rect 532 64274 604 64326
rect 656 64274 728 64326
rect 780 64274 929 64326
rect 71 64202 929 64274
rect 71 64150 232 64202
rect 284 64150 356 64202
rect 408 64150 480 64202
rect 532 64150 604 64202
rect 656 64150 728 64202
rect 780 64150 929 64202
rect 71 64078 929 64150
rect 71 64026 232 64078
rect 284 64026 356 64078
rect 408 64026 480 64078
rect 532 64026 604 64078
rect 656 64026 728 64078
rect 780 64026 929 64078
rect 71 63954 929 64026
rect 71 63902 232 63954
rect 284 63902 356 63954
rect 408 63902 480 63954
rect 532 63902 604 63954
rect 656 63902 728 63954
rect 780 63902 929 63954
rect 71 63830 929 63902
rect 71 63778 232 63830
rect 284 63778 356 63830
rect 408 63778 480 63830
rect 532 63778 604 63830
rect 656 63778 728 63830
rect 780 63778 929 63830
rect 71 63646 929 63778
rect 71 50548 82 63646
rect 918 50548 929 63646
rect 71 50416 929 50548
rect 71 50364 224 50416
rect 276 50364 348 50416
rect 400 50364 472 50416
rect 524 50364 596 50416
rect 648 50364 720 50416
rect 772 50364 929 50416
rect 71 50292 929 50364
rect 71 50240 224 50292
rect 276 50240 348 50292
rect 400 50240 472 50292
rect 524 50240 596 50292
rect 648 50240 720 50292
rect 772 50240 929 50292
rect 71 50168 929 50240
rect 71 50116 224 50168
rect 276 50116 348 50168
rect 400 50116 472 50168
rect 524 50116 596 50168
rect 648 50116 720 50168
rect 772 50116 929 50168
rect 71 50044 929 50116
rect 71 49992 224 50044
rect 276 49992 348 50044
rect 400 49992 472 50044
rect 524 49992 596 50044
rect 648 49992 720 50044
rect 772 49992 929 50044
rect 71 49920 929 49992
rect 71 49868 224 49920
rect 276 49868 348 49920
rect 400 49868 472 49920
rect 524 49868 596 49920
rect 648 49868 720 49920
rect 772 49868 929 49920
rect 71 49796 929 49868
rect 71 49744 224 49796
rect 276 49744 348 49796
rect 400 49744 472 49796
rect 524 49744 596 49796
rect 648 49744 720 49796
rect 772 49744 929 49796
rect 71 49672 929 49744
rect 71 49620 224 49672
rect 276 49620 348 49672
rect 400 49620 472 49672
rect 524 49620 596 49672
rect 648 49620 720 49672
rect 772 49620 929 49672
rect 71 49548 929 49620
rect 71 49496 224 49548
rect 276 49496 348 49548
rect 400 49496 472 49548
rect 524 49496 596 49548
rect 648 49496 720 49548
rect 772 49496 929 49548
rect 71 49424 929 49496
rect 71 49372 224 49424
rect 276 49372 348 49424
rect 400 49372 472 49424
rect 524 49372 596 49424
rect 648 49372 720 49424
rect 772 49372 929 49424
rect 71 49240 929 49372
rect 71 13276 82 49240
rect 918 13276 929 49240
rect 71 13265 929 13276
rect 71 13151 178 13265
rect -32 13119 178 13151
rect 824 13151 929 13265
rect 975 13151 1032 69897
rect 824 13119 1032 13151
rect -32 13108 1032 13119
<< via1 >>
rect 232 64770 284 64822
rect 356 64770 408 64822
rect 480 64770 532 64822
rect 604 64770 656 64822
rect 728 64770 780 64822
rect 232 64646 284 64698
rect 356 64646 408 64698
rect 480 64646 532 64698
rect 604 64646 656 64698
rect 728 64646 780 64698
rect 232 64522 284 64574
rect 356 64522 408 64574
rect 480 64522 532 64574
rect 604 64522 656 64574
rect 728 64522 780 64574
rect 232 64398 284 64450
rect 356 64398 408 64450
rect 480 64398 532 64450
rect 604 64398 656 64450
rect 728 64398 780 64450
rect 232 64274 284 64326
rect 356 64274 408 64326
rect 480 64274 532 64326
rect 604 64274 656 64326
rect 728 64274 780 64326
rect 232 64150 284 64202
rect 356 64150 408 64202
rect 480 64150 532 64202
rect 604 64150 656 64202
rect 728 64150 780 64202
rect 232 64026 284 64078
rect 356 64026 408 64078
rect 480 64026 532 64078
rect 604 64026 656 64078
rect 728 64026 780 64078
rect 232 63902 284 63954
rect 356 63902 408 63954
rect 480 63902 532 63954
rect 604 63902 656 63954
rect 728 63902 780 63954
rect 232 63778 284 63830
rect 356 63778 408 63830
rect 480 63778 532 63830
rect 604 63778 656 63830
rect 728 63778 780 63830
rect 224 50364 276 50416
rect 348 50364 400 50416
rect 472 50364 524 50416
rect 596 50364 648 50416
rect 720 50364 772 50416
rect 224 50240 276 50292
rect 348 50240 400 50292
rect 472 50240 524 50292
rect 596 50240 648 50292
rect 720 50240 772 50292
rect 224 50116 276 50168
rect 348 50116 400 50168
rect 472 50116 524 50168
rect 596 50116 648 50168
rect 720 50116 772 50168
rect 224 49992 276 50044
rect 348 49992 400 50044
rect 472 49992 524 50044
rect 596 49992 648 50044
rect 720 49992 772 50044
rect 224 49868 276 49920
rect 348 49868 400 49920
rect 472 49868 524 49920
rect 596 49868 648 49920
rect 720 49868 772 49920
rect 224 49744 276 49796
rect 348 49744 400 49796
rect 472 49744 524 49796
rect 596 49744 648 49796
rect 720 49744 772 49796
rect 224 49620 276 49672
rect 348 49620 400 49672
rect 472 49620 524 49672
rect 596 49620 648 49672
rect 720 49620 772 49672
rect 224 49496 276 49548
rect 348 49496 400 49548
rect 472 49496 524 49548
rect 596 49496 648 49548
rect 720 49496 772 49548
rect 224 49372 276 49424
rect 348 49372 400 49424
rect 472 49372 524 49424
rect 596 49372 648 49424
rect 720 49372 772 49424
<< metal2 >>
rect 0 64824 1000 65000
rect 0 64768 230 64824
rect 286 64768 354 64824
rect 410 64768 478 64824
rect 534 64768 602 64824
rect 658 64768 726 64824
rect 782 64768 1000 64824
rect 0 64700 1000 64768
rect 0 64644 230 64700
rect 286 64644 354 64700
rect 410 64644 478 64700
rect 534 64644 602 64700
rect 658 64644 726 64700
rect 782 64644 1000 64700
rect 0 64576 1000 64644
rect 0 64520 230 64576
rect 286 64520 354 64576
rect 410 64520 478 64576
rect 534 64520 602 64576
rect 658 64520 726 64576
rect 782 64520 1000 64576
rect 0 64452 1000 64520
rect 0 64396 230 64452
rect 286 64396 354 64452
rect 410 64396 478 64452
rect 534 64396 602 64452
rect 658 64396 726 64452
rect 782 64396 1000 64452
rect 0 64328 1000 64396
rect 0 64272 230 64328
rect 286 64272 354 64328
rect 410 64272 478 64328
rect 534 64272 602 64328
rect 658 64272 726 64328
rect 782 64272 1000 64328
rect 0 64204 1000 64272
rect 0 64148 230 64204
rect 286 64148 354 64204
rect 410 64148 478 64204
rect 534 64148 602 64204
rect 658 64148 726 64204
rect 782 64148 1000 64204
rect 0 64080 1000 64148
rect 0 64024 230 64080
rect 286 64024 354 64080
rect 410 64024 478 64080
rect 534 64024 602 64080
rect 658 64024 726 64080
rect 782 64024 1000 64080
rect 0 63956 1000 64024
rect 0 63900 230 63956
rect 286 63900 354 63956
rect 410 63900 478 63956
rect 534 63900 602 63956
rect 658 63900 726 63956
rect 782 63900 1000 63956
rect 0 63832 1000 63900
rect 0 63776 230 63832
rect 286 63776 354 63832
rect 410 63776 478 63832
rect 534 63776 602 63832
rect 658 63776 726 63832
rect 782 63776 1000 63832
rect 0 63600 1000 63776
rect 0 50418 1000 50600
rect 0 50362 222 50418
rect 278 50362 346 50418
rect 402 50362 470 50418
rect 526 50362 594 50418
rect 650 50362 718 50418
rect 774 50362 1000 50418
rect 0 50294 1000 50362
rect 0 50238 222 50294
rect 278 50238 346 50294
rect 402 50238 470 50294
rect 526 50238 594 50294
rect 650 50238 718 50294
rect 774 50238 1000 50294
rect 0 50170 1000 50238
rect 0 50114 222 50170
rect 278 50114 346 50170
rect 402 50114 470 50170
rect 526 50114 594 50170
rect 650 50114 718 50170
rect 774 50114 1000 50170
rect 0 50046 1000 50114
rect 0 49990 222 50046
rect 278 49990 346 50046
rect 402 49990 470 50046
rect 526 49990 594 50046
rect 650 49990 718 50046
rect 774 49990 1000 50046
rect 0 49922 1000 49990
rect 0 49866 222 49922
rect 278 49866 346 49922
rect 402 49866 470 49922
rect 526 49866 594 49922
rect 650 49866 718 49922
rect 774 49866 1000 49922
rect 0 49798 1000 49866
rect 0 49742 222 49798
rect 278 49742 346 49798
rect 402 49742 470 49798
rect 526 49742 594 49798
rect 650 49742 718 49798
rect 774 49742 1000 49798
rect 0 49674 1000 49742
rect 0 49618 222 49674
rect 278 49618 346 49674
rect 402 49618 470 49674
rect 526 49618 594 49674
rect 650 49618 718 49674
rect 774 49618 1000 49674
rect 0 49550 1000 49618
rect 0 49494 222 49550
rect 278 49494 346 49550
rect 402 49494 470 49550
rect 526 49494 594 49550
rect 650 49494 718 49550
rect 774 49494 1000 49550
rect 0 49426 1000 49494
rect 0 49370 222 49426
rect 278 49370 346 49426
rect 402 49370 470 49426
rect 526 49370 594 49426
rect 650 49370 718 49426
rect 774 49370 1000 49426
rect 0 49200 1000 49370
<< via2 >>
rect 230 64822 286 64824
rect 230 64770 232 64822
rect 232 64770 284 64822
rect 284 64770 286 64822
rect 230 64768 286 64770
rect 354 64822 410 64824
rect 354 64770 356 64822
rect 356 64770 408 64822
rect 408 64770 410 64822
rect 354 64768 410 64770
rect 478 64822 534 64824
rect 478 64770 480 64822
rect 480 64770 532 64822
rect 532 64770 534 64822
rect 478 64768 534 64770
rect 602 64822 658 64824
rect 602 64770 604 64822
rect 604 64770 656 64822
rect 656 64770 658 64822
rect 602 64768 658 64770
rect 726 64822 782 64824
rect 726 64770 728 64822
rect 728 64770 780 64822
rect 780 64770 782 64822
rect 726 64768 782 64770
rect 230 64698 286 64700
rect 230 64646 232 64698
rect 232 64646 284 64698
rect 284 64646 286 64698
rect 230 64644 286 64646
rect 354 64698 410 64700
rect 354 64646 356 64698
rect 356 64646 408 64698
rect 408 64646 410 64698
rect 354 64644 410 64646
rect 478 64698 534 64700
rect 478 64646 480 64698
rect 480 64646 532 64698
rect 532 64646 534 64698
rect 478 64644 534 64646
rect 602 64698 658 64700
rect 602 64646 604 64698
rect 604 64646 656 64698
rect 656 64646 658 64698
rect 602 64644 658 64646
rect 726 64698 782 64700
rect 726 64646 728 64698
rect 728 64646 780 64698
rect 780 64646 782 64698
rect 726 64644 782 64646
rect 230 64574 286 64576
rect 230 64522 232 64574
rect 232 64522 284 64574
rect 284 64522 286 64574
rect 230 64520 286 64522
rect 354 64574 410 64576
rect 354 64522 356 64574
rect 356 64522 408 64574
rect 408 64522 410 64574
rect 354 64520 410 64522
rect 478 64574 534 64576
rect 478 64522 480 64574
rect 480 64522 532 64574
rect 532 64522 534 64574
rect 478 64520 534 64522
rect 602 64574 658 64576
rect 602 64522 604 64574
rect 604 64522 656 64574
rect 656 64522 658 64574
rect 602 64520 658 64522
rect 726 64574 782 64576
rect 726 64522 728 64574
rect 728 64522 780 64574
rect 780 64522 782 64574
rect 726 64520 782 64522
rect 230 64450 286 64452
rect 230 64398 232 64450
rect 232 64398 284 64450
rect 284 64398 286 64450
rect 230 64396 286 64398
rect 354 64450 410 64452
rect 354 64398 356 64450
rect 356 64398 408 64450
rect 408 64398 410 64450
rect 354 64396 410 64398
rect 478 64450 534 64452
rect 478 64398 480 64450
rect 480 64398 532 64450
rect 532 64398 534 64450
rect 478 64396 534 64398
rect 602 64450 658 64452
rect 602 64398 604 64450
rect 604 64398 656 64450
rect 656 64398 658 64450
rect 602 64396 658 64398
rect 726 64450 782 64452
rect 726 64398 728 64450
rect 728 64398 780 64450
rect 780 64398 782 64450
rect 726 64396 782 64398
rect 230 64326 286 64328
rect 230 64274 232 64326
rect 232 64274 284 64326
rect 284 64274 286 64326
rect 230 64272 286 64274
rect 354 64326 410 64328
rect 354 64274 356 64326
rect 356 64274 408 64326
rect 408 64274 410 64326
rect 354 64272 410 64274
rect 478 64326 534 64328
rect 478 64274 480 64326
rect 480 64274 532 64326
rect 532 64274 534 64326
rect 478 64272 534 64274
rect 602 64326 658 64328
rect 602 64274 604 64326
rect 604 64274 656 64326
rect 656 64274 658 64326
rect 602 64272 658 64274
rect 726 64326 782 64328
rect 726 64274 728 64326
rect 728 64274 780 64326
rect 780 64274 782 64326
rect 726 64272 782 64274
rect 230 64202 286 64204
rect 230 64150 232 64202
rect 232 64150 284 64202
rect 284 64150 286 64202
rect 230 64148 286 64150
rect 354 64202 410 64204
rect 354 64150 356 64202
rect 356 64150 408 64202
rect 408 64150 410 64202
rect 354 64148 410 64150
rect 478 64202 534 64204
rect 478 64150 480 64202
rect 480 64150 532 64202
rect 532 64150 534 64202
rect 478 64148 534 64150
rect 602 64202 658 64204
rect 602 64150 604 64202
rect 604 64150 656 64202
rect 656 64150 658 64202
rect 602 64148 658 64150
rect 726 64202 782 64204
rect 726 64150 728 64202
rect 728 64150 780 64202
rect 780 64150 782 64202
rect 726 64148 782 64150
rect 230 64078 286 64080
rect 230 64026 232 64078
rect 232 64026 284 64078
rect 284 64026 286 64078
rect 230 64024 286 64026
rect 354 64078 410 64080
rect 354 64026 356 64078
rect 356 64026 408 64078
rect 408 64026 410 64078
rect 354 64024 410 64026
rect 478 64078 534 64080
rect 478 64026 480 64078
rect 480 64026 532 64078
rect 532 64026 534 64078
rect 478 64024 534 64026
rect 602 64078 658 64080
rect 602 64026 604 64078
rect 604 64026 656 64078
rect 656 64026 658 64078
rect 602 64024 658 64026
rect 726 64078 782 64080
rect 726 64026 728 64078
rect 728 64026 780 64078
rect 780 64026 782 64078
rect 726 64024 782 64026
rect 230 63954 286 63956
rect 230 63902 232 63954
rect 232 63902 284 63954
rect 284 63902 286 63954
rect 230 63900 286 63902
rect 354 63954 410 63956
rect 354 63902 356 63954
rect 356 63902 408 63954
rect 408 63902 410 63954
rect 354 63900 410 63902
rect 478 63954 534 63956
rect 478 63902 480 63954
rect 480 63902 532 63954
rect 532 63902 534 63954
rect 478 63900 534 63902
rect 602 63954 658 63956
rect 602 63902 604 63954
rect 604 63902 656 63954
rect 656 63902 658 63954
rect 602 63900 658 63902
rect 726 63954 782 63956
rect 726 63902 728 63954
rect 728 63902 780 63954
rect 780 63902 782 63954
rect 726 63900 782 63902
rect 230 63830 286 63832
rect 230 63778 232 63830
rect 232 63778 284 63830
rect 284 63778 286 63830
rect 230 63776 286 63778
rect 354 63830 410 63832
rect 354 63778 356 63830
rect 356 63778 408 63830
rect 408 63778 410 63830
rect 354 63776 410 63778
rect 478 63830 534 63832
rect 478 63778 480 63830
rect 480 63778 532 63830
rect 532 63778 534 63830
rect 478 63776 534 63778
rect 602 63830 658 63832
rect 602 63778 604 63830
rect 604 63778 656 63830
rect 656 63778 658 63830
rect 602 63776 658 63778
rect 726 63830 782 63832
rect 726 63778 728 63830
rect 728 63778 780 63830
rect 780 63778 782 63830
rect 726 63776 782 63778
rect 222 50416 278 50418
rect 222 50364 224 50416
rect 224 50364 276 50416
rect 276 50364 278 50416
rect 222 50362 278 50364
rect 346 50416 402 50418
rect 346 50364 348 50416
rect 348 50364 400 50416
rect 400 50364 402 50416
rect 346 50362 402 50364
rect 470 50416 526 50418
rect 470 50364 472 50416
rect 472 50364 524 50416
rect 524 50364 526 50416
rect 470 50362 526 50364
rect 594 50416 650 50418
rect 594 50364 596 50416
rect 596 50364 648 50416
rect 648 50364 650 50416
rect 594 50362 650 50364
rect 718 50416 774 50418
rect 718 50364 720 50416
rect 720 50364 772 50416
rect 772 50364 774 50416
rect 718 50362 774 50364
rect 222 50292 278 50294
rect 222 50240 224 50292
rect 224 50240 276 50292
rect 276 50240 278 50292
rect 222 50238 278 50240
rect 346 50292 402 50294
rect 346 50240 348 50292
rect 348 50240 400 50292
rect 400 50240 402 50292
rect 346 50238 402 50240
rect 470 50292 526 50294
rect 470 50240 472 50292
rect 472 50240 524 50292
rect 524 50240 526 50292
rect 470 50238 526 50240
rect 594 50292 650 50294
rect 594 50240 596 50292
rect 596 50240 648 50292
rect 648 50240 650 50292
rect 594 50238 650 50240
rect 718 50292 774 50294
rect 718 50240 720 50292
rect 720 50240 772 50292
rect 772 50240 774 50292
rect 718 50238 774 50240
rect 222 50168 278 50170
rect 222 50116 224 50168
rect 224 50116 276 50168
rect 276 50116 278 50168
rect 222 50114 278 50116
rect 346 50168 402 50170
rect 346 50116 348 50168
rect 348 50116 400 50168
rect 400 50116 402 50168
rect 346 50114 402 50116
rect 470 50168 526 50170
rect 470 50116 472 50168
rect 472 50116 524 50168
rect 524 50116 526 50168
rect 470 50114 526 50116
rect 594 50168 650 50170
rect 594 50116 596 50168
rect 596 50116 648 50168
rect 648 50116 650 50168
rect 594 50114 650 50116
rect 718 50168 774 50170
rect 718 50116 720 50168
rect 720 50116 772 50168
rect 772 50116 774 50168
rect 718 50114 774 50116
rect 222 50044 278 50046
rect 222 49992 224 50044
rect 224 49992 276 50044
rect 276 49992 278 50044
rect 222 49990 278 49992
rect 346 50044 402 50046
rect 346 49992 348 50044
rect 348 49992 400 50044
rect 400 49992 402 50044
rect 346 49990 402 49992
rect 470 50044 526 50046
rect 470 49992 472 50044
rect 472 49992 524 50044
rect 524 49992 526 50044
rect 470 49990 526 49992
rect 594 50044 650 50046
rect 594 49992 596 50044
rect 596 49992 648 50044
rect 648 49992 650 50044
rect 594 49990 650 49992
rect 718 50044 774 50046
rect 718 49992 720 50044
rect 720 49992 772 50044
rect 772 49992 774 50044
rect 718 49990 774 49992
rect 222 49920 278 49922
rect 222 49868 224 49920
rect 224 49868 276 49920
rect 276 49868 278 49920
rect 222 49866 278 49868
rect 346 49920 402 49922
rect 346 49868 348 49920
rect 348 49868 400 49920
rect 400 49868 402 49920
rect 346 49866 402 49868
rect 470 49920 526 49922
rect 470 49868 472 49920
rect 472 49868 524 49920
rect 524 49868 526 49920
rect 470 49866 526 49868
rect 594 49920 650 49922
rect 594 49868 596 49920
rect 596 49868 648 49920
rect 648 49868 650 49920
rect 594 49866 650 49868
rect 718 49920 774 49922
rect 718 49868 720 49920
rect 720 49868 772 49920
rect 772 49868 774 49920
rect 718 49866 774 49868
rect 222 49796 278 49798
rect 222 49744 224 49796
rect 224 49744 276 49796
rect 276 49744 278 49796
rect 222 49742 278 49744
rect 346 49796 402 49798
rect 346 49744 348 49796
rect 348 49744 400 49796
rect 400 49744 402 49796
rect 346 49742 402 49744
rect 470 49796 526 49798
rect 470 49744 472 49796
rect 472 49744 524 49796
rect 524 49744 526 49796
rect 470 49742 526 49744
rect 594 49796 650 49798
rect 594 49744 596 49796
rect 596 49744 648 49796
rect 648 49744 650 49796
rect 594 49742 650 49744
rect 718 49796 774 49798
rect 718 49744 720 49796
rect 720 49744 772 49796
rect 772 49744 774 49796
rect 718 49742 774 49744
rect 222 49672 278 49674
rect 222 49620 224 49672
rect 224 49620 276 49672
rect 276 49620 278 49672
rect 222 49618 278 49620
rect 346 49672 402 49674
rect 346 49620 348 49672
rect 348 49620 400 49672
rect 400 49620 402 49672
rect 346 49618 402 49620
rect 470 49672 526 49674
rect 470 49620 472 49672
rect 472 49620 524 49672
rect 524 49620 526 49672
rect 470 49618 526 49620
rect 594 49672 650 49674
rect 594 49620 596 49672
rect 596 49620 648 49672
rect 648 49620 650 49672
rect 594 49618 650 49620
rect 718 49672 774 49674
rect 718 49620 720 49672
rect 720 49620 772 49672
rect 772 49620 774 49672
rect 718 49618 774 49620
rect 222 49548 278 49550
rect 222 49496 224 49548
rect 224 49496 276 49548
rect 276 49496 278 49548
rect 222 49494 278 49496
rect 346 49548 402 49550
rect 346 49496 348 49548
rect 348 49496 400 49548
rect 400 49496 402 49548
rect 346 49494 402 49496
rect 470 49548 526 49550
rect 470 49496 472 49548
rect 472 49496 524 49548
rect 524 49496 526 49548
rect 470 49494 526 49496
rect 594 49548 650 49550
rect 594 49496 596 49548
rect 596 49496 648 49548
rect 648 49496 650 49548
rect 594 49494 650 49496
rect 718 49548 774 49550
rect 718 49496 720 49548
rect 720 49496 772 49548
rect 772 49496 774 49548
rect 718 49494 774 49496
rect 222 49424 278 49426
rect 222 49372 224 49424
rect 224 49372 276 49424
rect 276 49372 278 49424
rect 222 49370 278 49372
rect 346 49424 402 49426
rect 346 49372 348 49424
rect 348 49372 400 49424
rect 400 49372 402 49424
rect 346 49370 402 49372
rect 470 49424 526 49426
rect 470 49372 472 49424
rect 472 49372 524 49424
rect 524 49372 526 49424
rect 470 49370 526 49372
rect 594 49424 650 49426
rect 594 49372 596 49424
rect 596 49372 648 49424
rect 648 49372 650 49424
rect 594 49370 650 49372
rect 718 49424 774 49426
rect 718 49372 720 49424
rect 720 49372 772 49424
rect 772 49372 774 49424
rect 718 49370 774 49372
<< metal3 >>
rect 0 64824 1000 65000
rect 0 64768 230 64824
rect 286 64768 354 64824
rect 410 64768 478 64824
rect 534 64768 602 64824
rect 658 64768 726 64824
rect 782 64768 1000 64824
rect 0 64700 1000 64768
rect 0 64644 230 64700
rect 286 64644 354 64700
rect 410 64644 478 64700
rect 534 64644 602 64700
rect 658 64644 726 64700
rect 782 64644 1000 64700
rect 0 64576 1000 64644
rect 0 64520 230 64576
rect 286 64520 354 64576
rect 410 64520 478 64576
rect 534 64520 602 64576
rect 658 64520 726 64576
rect 782 64520 1000 64576
rect 0 64452 1000 64520
rect 0 64396 230 64452
rect 286 64396 354 64452
rect 410 64396 478 64452
rect 534 64396 602 64452
rect 658 64396 726 64452
rect 782 64396 1000 64452
rect 0 64328 1000 64396
rect 0 64272 230 64328
rect 286 64272 354 64328
rect 410 64272 478 64328
rect 534 64272 602 64328
rect 658 64272 726 64328
rect 782 64272 1000 64328
rect 0 64204 1000 64272
rect 0 64148 230 64204
rect 286 64148 354 64204
rect 410 64148 478 64204
rect 534 64148 602 64204
rect 658 64148 726 64204
rect 782 64148 1000 64204
rect 0 64080 1000 64148
rect 0 64024 230 64080
rect 286 64024 354 64080
rect 410 64024 478 64080
rect 534 64024 602 64080
rect 658 64024 726 64080
rect 782 64024 1000 64080
rect 0 63956 1000 64024
rect 0 63900 230 63956
rect 286 63900 354 63956
rect 410 63900 478 63956
rect 534 63900 602 63956
rect 658 63900 726 63956
rect 782 63900 1000 63956
rect 0 63832 1000 63900
rect 0 63776 230 63832
rect 286 63776 354 63832
rect 410 63776 478 63832
rect 534 63776 602 63832
rect 658 63776 726 63832
rect 782 63776 1000 63832
rect 0 63600 1000 63776
rect 0 50418 1000 50600
rect 0 50362 222 50418
rect 278 50362 346 50418
rect 402 50362 470 50418
rect 526 50362 594 50418
rect 650 50362 718 50418
rect 774 50362 1000 50418
rect 0 50294 1000 50362
rect 0 50238 222 50294
rect 278 50238 346 50294
rect 402 50238 470 50294
rect 526 50238 594 50294
rect 650 50238 718 50294
rect 774 50238 1000 50294
rect 0 50170 1000 50238
rect 0 50114 222 50170
rect 278 50114 346 50170
rect 402 50114 470 50170
rect 526 50114 594 50170
rect 650 50114 718 50170
rect 774 50114 1000 50170
rect 0 50046 1000 50114
rect 0 49990 222 50046
rect 278 49990 346 50046
rect 402 49990 470 50046
rect 526 49990 594 50046
rect 650 49990 718 50046
rect 774 49990 1000 50046
rect 0 49922 1000 49990
rect 0 49866 222 49922
rect 278 49866 346 49922
rect 402 49866 470 49922
rect 526 49866 594 49922
rect 650 49866 718 49922
rect 774 49866 1000 49922
rect 0 49798 1000 49866
rect 0 49742 222 49798
rect 278 49742 346 49798
rect 402 49742 470 49798
rect 526 49742 594 49798
rect 650 49742 718 49798
rect 774 49742 1000 49798
rect 0 49674 1000 49742
rect 0 49618 222 49674
rect 278 49618 346 49674
rect 402 49618 470 49674
rect 526 49618 594 49674
rect 650 49618 718 49674
rect 774 49618 1000 49674
rect 0 49550 1000 49618
rect 0 49494 222 49550
rect 278 49494 346 49550
rect 402 49494 470 49550
rect 526 49494 594 49550
rect 650 49494 718 49550
rect 774 49494 1000 49550
rect 0 49426 1000 49494
rect 0 49370 222 49426
rect 278 49370 346 49426
rect 402 49370 470 49426
rect 526 49370 594 49426
rect 650 49370 718 49426
rect 774 49370 1000 49426
rect 0 49200 1000 49370
use M1_PSUB_CDNS_406619531455  M1_PSUB_CDNS_406619531455_0
timestamp 1755724134
transform -1 0 48 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_406619531455  M1_PSUB_CDNS_406619531455_1
timestamp 1755724134
transform 1 0 952 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_4066195314516  M1_PSUB_CDNS_4066195314516_0
timestamp 1755724134
transform 1 0 501 0 -1 13192
box 0 0 1 1
use M1_PSUB_CDNS_4066195314516  M1_PSUB_CDNS_4066195314516_1
timestamp 1755724134
transform 1 0 501 0 1 69873
box 0 0 1 1
use M2_M1_CDNS_4066195314542  M2_M1_CDNS_4066195314542_0
timestamp 1755724134
transform 1 0 498 0 1 49894
box 0 0 1 1
use M2_M1_CDNS_4066195314542  M2_M1_CDNS_4066195314542_1
timestamp 1755724134
transform 1 0 506 0 1 64300
box 0 0 1 1
use M3_M2_CDNS_4066195314543  M3_M2_CDNS_4066195314543_0
timestamp 1755724134
transform 1 0 498 0 1 49894
box 0 0 1 1
use M3_M2_CDNS_4066195314543  M3_M2_CDNS_4066195314543_1
timestamp 1755724134
transform 1 0 506 0 1 64300
box 0 0 1 1
use POLY_SUB_FILL_3  POLY_SUB_FILL_3_0
array 0 0 0 0 96 574
timestamp 1755724134
transform 1 0 187 0 1 13813
box -127 -235 772 615
<< labels >>
rlabel metal3 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 510 50023 510 50023 4 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string GDS_END 3665576
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3663940
<< end >>
