magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 4342 870
<< pwell >>
rect -86 -86 4342 352
<< mvnmos >>
rect 124 155 244 228
rect 348 155 468 228
rect 572 155 692 228
rect 796 155 916 228
rect 1020 155 1140 228
rect 1504 132 1624 228
rect 1728 132 1848 228
rect 1952 132 2072 228
rect 2176 132 2296 228
rect 2400 132 2520 228
rect 2624 132 2744 228
rect 2848 132 2968 228
rect 3072 132 3192 228
rect 3296 132 3416 228
rect 3520 132 3640 228
rect 3744 132 3864 228
rect 3968 132 4088 228
<< mvpmos >>
rect 124 552 224 716
rect 348 552 448 716
rect 572 552 672 716
rect 796 552 896 716
rect 1020 552 1120 716
rect 1244 552 1344 716
rect 1504 472 1604 716
rect 1728 472 1828 716
rect 1952 472 2052 716
rect 2176 472 2276 716
rect 2400 472 2500 716
rect 2624 472 2724 716
rect 2848 472 2948 716
rect 3072 472 3172 716
rect 3296 472 3396 716
rect 3520 472 3620 716
rect 3744 472 3844 716
rect 3968 472 4068 716
<< mvndiff >>
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 155 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 155 348 169
rect 468 215 572 228
rect 468 169 497 215
rect 543 169 572 215
rect 468 155 572 169
rect 692 215 796 228
rect 692 169 721 215
rect 767 169 796 215
rect 692 155 796 169
rect 916 215 1020 228
rect 916 169 945 215
rect 991 169 1020 215
rect 916 155 1020 169
rect 1140 215 1228 228
rect 1140 169 1169 215
rect 1215 169 1228 215
rect 1140 155 1228 169
rect 1416 215 1504 228
rect 1416 169 1429 215
rect 1475 169 1504 215
rect 1416 132 1504 169
rect 1624 197 1728 228
rect 1624 151 1653 197
rect 1699 151 1728 197
rect 1624 132 1728 151
rect 1848 197 1952 228
rect 1848 151 1877 197
rect 1923 151 1952 197
rect 1848 132 1952 151
rect 2072 197 2176 228
rect 2072 151 2101 197
rect 2147 151 2176 197
rect 2072 132 2176 151
rect 2296 197 2400 228
rect 2296 151 2325 197
rect 2371 151 2400 197
rect 2296 132 2400 151
rect 2520 197 2624 228
rect 2520 151 2549 197
rect 2595 151 2624 197
rect 2520 132 2624 151
rect 2744 197 2848 228
rect 2744 151 2773 197
rect 2819 151 2848 197
rect 2744 132 2848 151
rect 2968 197 3072 228
rect 2968 151 2997 197
rect 3043 151 3072 197
rect 2968 132 3072 151
rect 3192 197 3296 228
rect 3192 151 3221 197
rect 3267 151 3296 197
rect 3192 132 3296 151
rect 3416 197 3520 228
rect 3416 151 3445 197
rect 3491 151 3520 197
rect 3416 132 3520 151
rect 3640 197 3744 228
rect 3640 151 3669 197
rect 3715 151 3744 197
rect 3640 132 3744 151
rect 3864 197 3968 228
rect 3864 151 3893 197
rect 3939 151 3968 197
rect 3864 132 3968 151
rect 4088 197 4176 228
rect 4088 151 4117 197
rect 4163 151 4176 197
rect 4088 132 4176 151
<< mvpdiff >>
rect 36 703 124 716
rect 36 657 49 703
rect 95 657 124 703
rect 36 552 124 657
rect 224 665 348 716
rect 224 619 253 665
rect 299 619 348 665
rect 224 552 348 619
rect 448 667 572 716
rect 448 621 477 667
rect 523 621 572 667
rect 448 552 572 621
rect 672 665 796 716
rect 672 619 701 665
rect 747 619 796 665
rect 672 552 796 619
rect 896 667 1020 716
rect 896 621 925 667
rect 971 621 1020 667
rect 896 552 1020 621
rect 1120 665 1244 716
rect 1120 619 1149 665
rect 1195 619 1244 665
rect 1120 552 1244 619
rect 1344 703 1504 716
rect 1344 657 1429 703
rect 1475 657 1504 703
rect 1344 552 1504 657
rect 1424 472 1504 552
rect 1604 665 1728 716
rect 1604 525 1653 665
rect 1699 525 1728 665
rect 1604 472 1728 525
rect 1828 703 1952 716
rect 1828 657 1857 703
rect 1903 657 1952 703
rect 1828 472 1952 657
rect 2052 665 2176 716
rect 2052 525 2081 665
rect 2127 525 2176 665
rect 2052 472 2176 525
rect 2276 703 2400 716
rect 2276 657 2305 703
rect 2351 657 2400 703
rect 2276 472 2400 657
rect 2500 665 2624 716
rect 2500 525 2529 665
rect 2575 525 2624 665
rect 2500 472 2624 525
rect 2724 703 2848 716
rect 2724 657 2753 703
rect 2799 657 2848 703
rect 2724 472 2848 657
rect 2948 665 3072 716
rect 2948 525 2977 665
rect 3023 525 3072 665
rect 2948 472 3072 525
rect 3172 703 3296 716
rect 3172 657 3201 703
rect 3247 657 3296 703
rect 3172 472 3296 657
rect 3396 665 3520 716
rect 3396 525 3425 665
rect 3471 525 3520 665
rect 3396 472 3520 525
rect 3620 703 3744 716
rect 3620 657 3649 703
rect 3695 657 3744 703
rect 3620 472 3744 657
rect 3844 665 3968 716
rect 3844 525 3873 665
rect 3919 525 3968 665
rect 3844 472 3968 525
rect 4068 703 4156 716
rect 4068 563 4097 703
rect 4143 563 4156 703
rect 4068 472 4156 563
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 497 169 543 215
rect 721 169 767 215
rect 945 169 991 215
rect 1169 169 1215 215
rect 1429 169 1475 215
rect 1653 151 1699 197
rect 1877 151 1923 197
rect 2101 151 2147 197
rect 2325 151 2371 197
rect 2549 151 2595 197
rect 2773 151 2819 197
rect 2997 151 3043 197
rect 3221 151 3267 197
rect 3445 151 3491 197
rect 3669 151 3715 197
rect 3893 151 3939 197
rect 4117 151 4163 197
<< mvpdiffc >>
rect 49 657 95 703
rect 253 619 299 665
rect 477 621 523 667
rect 701 619 747 665
rect 925 621 971 667
rect 1149 619 1195 665
rect 1429 657 1475 703
rect 1653 525 1699 665
rect 1857 657 1903 703
rect 2081 525 2127 665
rect 2305 657 2351 703
rect 2529 525 2575 665
rect 2753 657 2799 703
rect 2977 525 3023 665
rect 3201 657 3247 703
rect 3425 525 3471 665
rect 3649 657 3695 703
rect 3873 525 3919 665
rect 4097 563 4143 703
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1504 716 1604 760
rect 1728 716 1828 760
rect 1952 716 2052 760
rect 2176 716 2276 760
rect 2400 716 2500 760
rect 2624 716 2724 760
rect 2848 716 2948 760
rect 3072 716 3172 760
rect 3296 716 3396 760
rect 3520 716 3620 760
rect 3744 716 3844 760
rect 3968 716 4068 760
rect 124 412 224 552
rect 348 412 448 552
rect 572 412 672 552
rect 796 412 896 552
rect 1020 412 1120 552
rect 1244 412 1344 552
rect 124 399 1344 412
rect 124 353 181 399
rect 1167 353 1344 399
rect 124 340 1344 353
rect 1504 412 1604 472
rect 1728 412 1828 472
rect 1952 412 2052 472
rect 2176 412 2276 472
rect 2400 412 2500 472
rect 2624 412 2724 472
rect 2848 412 2948 472
rect 3072 412 3172 472
rect 3296 412 3396 472
rect 3520 412 3620 472
rect 3744 412 3844 472
rect 3968 412 4068 472
rect 1504 399 4088 412
rect 1504 353 1517 399
rect 2597 353 3089 399
rect 4075 353 4088 399
rect 1504 340 4088 353
rect 124 228 244 340
rect 348 228 468 340
rect 572 228 692 340
rect 796 228 916 340
rect 1020 228 1140 340
rect 1504 228 1624 340
rect 1728 228 1848 340
rect 1952 228 2072 340
rect 2176 228 2296 340
rect 2400 228 2520 340
rect 2624 228 2744 340
rect 2848 228 2968 340
rect 3072 228 3192 340
rect 3296 228 3416 340
rect 3520 228 3640 340
rect 3744 228 3864 340
rect 3968 228 4088 340
rect 124 94 244 155
rect 348 94 468 155
rect 572 94 692 155
rect 796 94 916 155
rect 1020 94 1140 155
rect 1504 88 1624 132
rect 1728 88 1848 132
rect 1952 88 2072 132
rect 2176 88 2296 132
rect 2400 88 2520 132
rect 2624 88 2744 132
rect 2848 88 2968 132
rect 3072 88 3192 132
rect 3296 88 3416 132
rect 3520 88 3640 132
rect 3744 88 3864 132
rect 3968 88 4088 132
<< polycontact >>
rect 181 353 1167 399
rect 1517 353 2597 399
rect 3089 353 4075 399
<< metal1 >>
rect 0 724 4256 844
rect 49 703 95 724
rect 49 646 95 657
rect 253 665 299 678
rect 253 552 299 619
rect 477 667 523 724
rect 477 610 523 621
rect 701 665 747 678
rect 701 552 747 619
rect 925 667 971 724
rect 1429 703 1475 724
rect 925 610 971 621
rect 1149 665 1195 678
rect 1857 703 1903 724
rect 1429 646 1475 657
rect 1653 665 1699 678
rect 1149 552 1195 619
rect 253 506 1319 552
rect 124 399 1214 430
rect 124 353 181 399
rect 1167 353 1214 399
rect 1273 413 1319 506
rect 2305 703 2351 724
rect 1857 646 1903 657
rect 2081 665 2127 678
rect 1699 525 2081 600
rect 2753 703 2799 724
rect 2305 646 2351 657
rect 2529 665 2575 678
rect 2127 525 2529 600
rect 3201 703 3247 724
rect 2753 646 2799 657
rect 2977 665 3023 678
rect 2575 525 2977 600
rect 3649 703 3695 724
rect 3201 646 3247 657
rect 3425 665 3471 678
rect 3023 525 3425 600
rect 4097 703 4143 724
rect 3649 646 3695 657
rect 3873 665 3919 678
rect 3471 525 3873 600
rect 4097 552 4143 563
rect 1653 499 3919 525
rect 1273 399 2618 413
rect 1273 353 1517 399
rect 2597 353 2618 399
rect 1273 307 1319 353
rect 2766 307 2946 499
rect 3078 399 4086 413
rect 3078 353 3089 399
rect 4075 353 4086 399
rect 262 261 1319 307
rect 262 215 330 261
rect 710 215 778 261
rect 1158 215 1226 261
rect 1653 243 3939 307
rect 38 169 49 215
rect 95 169 106 215
rect 262 169 273 215
rect 319 169 330 215
rect 486 169 497 215
rect 543 169 554 215
rect 710 169 721 215
rect 767 169 778 215
rect 934 169 945 215
rect 991 169 1002 215
rect 1158 169 1169 215
rect 1215 169 1226 215
rect 1418 169 1429 215
rect 1475 169 1486 215
rect 38 60 106 169
rect 486 60 554 169
rect 934 60 1002 169
rect 1418 60 1486 169
rect 1653 197 1699 243
rect 2101 197 2147 243
rect 2549 197 2595 243
rect 2997 197 3043 243
rect 3445 197 3491 243
rect 3893 197 3939 243
rect 1653 138 1699 151
rect 1866 151 1877 197
rect 1923 151 1934 197
rect 1866 60 1934 151
rect 2101 138 2147 151
rect 2314 151 2325 197
rect 2371 151 2382 197
rect 2314 60 2382 151
rect 2549 138 2595 151
rect 2762 151 2773 197
rect 2819 151 2830 197
rect 2762 60 2830 151
rect 2997 138 3043 151
rect 3210 151 3221 197
rect 3267 151 3278 197
rect 3210 60 3278 151
rect 3445 138 3491 151
rect 3658 151 3669 197
rect 3715 151 3726 197
rect 3658 60 3726 151
rect 3893 138 3939 151
rect 4106 151 4117 197
rect 4163 151 4174 197
rect 4106 60 4174 151
rect 0 -60 4256 60
<< labels >>
flabel metal1 s 0 724 4256 844 0 FreeSans 600 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 1418 197 1486 215 0 FreeSans 600 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3873 600 3919 678 0 FreeSans 600 0 0 0 Z
port 2 nsew default output
flabel metal1 s 124 353 1214 430 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 3425 600 3471 678 1 Z
port 2 nsew default output
rlabel metal1 s 2977 600 3023 678 1 Z
port 2 nsew default output
rlabel metal1 s 2529 600 2575 678 1 Z
port 2 nsew default output
rlabel metal1 s 2081 600 2127 678 1 Z
port 2 nsew default output
rlabel metal1 s 1653 600 1699 678 1 Z
port 2 nsew default output
rlabel metal1 s 1653 499 3919 600 1 Z
port 2 nsew default output
rlabel metal1 s 2766 307 2946 499 1 Z
port 2 nsew default output
rlabel metal1 s 1653 243 3939 307 1 Z
port 2 nsew default output
rlabel metal1 s 3893 138 3939 243 1 Z
port 2 nsew default output
rlabel metal1 s 3445 138 3491 243 1 Z
port 2 nsew default output
rlabel metal1 s 2997 138 3043 243 1 Z
port 2 nsew default output
rlabel metal1 s 2549 138 2595 243 1 Z
port 2 nsew default output
rlabel metal1 s 2101 138 2147 243 1 Z
port 2 nsew default output
rlabel metal1 s 1653 138 1699 243 1 Z
port 2 nsew default output
rlabel metal1 s 4097 646 4143 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3649 646 3695 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3201 646 3247 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2753 646 2799 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2305 646 2351 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1857 646 1903 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1429 646 1475 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4097 610 4143 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 610 971 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 610 523 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4097 552 4143 610 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 934 197 1002 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 197 554 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 197 106 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4106 60 4174 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3658 60 3726 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3210 60 3278 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2762 60 2830 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2314 60 2382 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1866 60 1934 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1418 60 1486 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string GDS_END 789406
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 780202
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
