magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 3782 870
<< pwell >>
rect -86 -86 3782 352
<< mvnmos >>
rect 124 90 244 232
rect 392 156 512 232
rect 560 156 680 232
rect 728 156 848 232
rect 952 156 1072 232
rect 1176 156 1296 232
rect 1488 156 1608 232
rect 1712 156 1832 232
rect 2080 156 2200 232
rect 2392 156 2512 232
rect 2704 156 2824 232
rect 2928 156 3048 232
rect 3096 156 3216 232
rect 3364 69 3484 232
<< mvpmos >>
rect 144 472 244 715
rect 412 496 512 628
rect 580 496 680 628
rect 748 496 848 628
rect 972 496 1072 628
rect 1196 496 1296 628
rect 1488 496 1588 628
rect 1692 496 1792 628
rect 2100 472 2200 612
rect 2392 472 2492 612
rect 2704 472 2804 612
rect 2928 472 3028 612
rect 3096 472 3196 612
rect 3364 472 3464 715
<< mvndiff >>
rect 36 218 124 232
rect 36 172 49 218
rect 95 172 124 218
rect 36 90 124 172
rect 244 163 392 232
rect 244 117 273 163
rect 319 156 392 163
rect 512 156 560 232
rect 680 156 728 232
rect 848 219 952 232
rect 848 173 877 219
rect 923 173 952 219
rect 848 156 952 173
rect 1072 219 1176 232
rect 1072 173 1101 219
rect 1147 173 1176 219
rect 1072 156 1176 173
rect 1296 183 1488 232
rect 1296 156 1369 183
rect 319 117 332 156
rect 244 90 332 117
rect 1356 137 1369 156
rect 1415 156 1488 183
rect 1608 219 1712 232
rect 1608 173 1637 219
rect 1683 173 1712 219
rect 1608 156 1712 173
rect 1832 218 1920 232
rect 1832 172 1861 218
rect 1907 172 1920 218
rect 1832 156 1920 172
rect 1992 215 2080 232
rect 1992 169 2005 215
rect 2051 169 2080 215
rect 1992 156 2080 169
rect 2200 183 2392 232
rect 2200 156 2273 183
rect 1415 137 1428 156
rect 1356 124 1428 137
rect 2260 137 2273 156
rect 2319 156 2392 183
rect 2512 183 2704 232
rect 2512 156 2585 183
rect 2319 137 2332 156
rect 2260 124 2332 137
rect 2572 137 2585 156
rect 2631 156 2704 183
rect 2824 215 2928 232
rect 2824 169 2853 215
rect 2899 169 2928 215
rect 2824 156 2928 169
rect 3048 156 3096 232
rect 3216 156 3364 232
rect 2631 137 2644 156
rect 2572 124 2644 137
rect 3276 142 3364 156
rect 3276 96 3289 142
rect 3335 96 3364 142
rect 3276 69 3364 96
rect 3484 215 3572 232
rect 3484 169 3513 215
rect 3559 169 3572 215
rect 3484 69 3572 169
<< mvpdiff >>
rect 56 663 144 715
rect 56 523 69 663
rect 115 523 144 663
rect 56 472 144 523
rect 244 689 332 715
rect 244 643 273 689
rect 319 643 332 689
rect 244 628 332 643
rect 1356 647 1428 660
rect 1356 628 1369 647
rect 244 496 412 628
rect 512 496 580 628
rect 680 496 748 628
rect 848 558 972 628
rect 848 512 877 558
rect 923 512 972 558
rect 848 496 972 512
rect 1072 558 1196 628
rect 1072 512 1121 558
rect 1167 512 1196 558
rect 1072 496 1196 512
rect 1296 601 1369 628
rect 1415 628 1428 647
rect 1415 601 1488 628
rect 1296 496 1488 601
rect 1588 558 1692 628
rect 1588 512 1617 558
rect 1663 512 1692 558
rect 1588 496 1692 512
rect 1792 598 1880 628
rect 2260 647 2332 660
rect 2260 612 2273 647
rect 1792 552 1821 598
rect 1867 552 1880 598
rect 1792 496 1880 552
rect 2012 555 2100 612
rect 2012 509 2025 555
rect 2071 509 2100 555
rect 244 472 324 496
rect 2012 472 2100 509
rect 2200 601 2273 612
rect 2319 612 2332 647
rect 3276 655 3364 715
rect 3276 612 3289 655
rect 2319 601 2392 612
rect 2200 472 2392 601
rect 2492 555 2704 612
rect 2492 509 2521 555
rect 2567 509 2629 555
rect 2675 509 2704 555
rect 2492 472 2704 509
rect 2804 534 2928 612
rect 2804 488 2833 534
rect 2879 488 2928 534
rect 2804 472 2928 488
rect 3028 472 3096 612
rect 3196 515 3289 612
rect 3335 515 3364 655
rect 3196 472 3364 515
rect 3464 655 3552 715
rect 3464 515 3493 655
rect 3539 515 3552 655
rect 3464 472 3552 515
<< mvndiffc >>
rect 49 172 95 218
rect 273 117 319 163
rect 877 173 923 219
rect 1101 173 1147 219
rect 1369 137 1415 183
rect 1637 173 1683 219
rect 1861 172 1907 218
rect 2005 169 2051 215
rect 2273 137 2319 183
rect 2585 137 2631 183
rect 2853 169 2899 215
rect 3289 96 3335 142
rect 3513 169 3559 215
<< mvpdiffc >>
rect 69 523 115 663
rect 273 643 319 689
rect 877 512 923 558
rect 1121 512 1167 558
rect 1369 601 1415 647
rect 1617 512 1663 558
rect 1821 552 1867 598
rect 2025 509 2071 555
rect 2273 601 2319 647
rect 2521 509 2567 555
rect 2629 509 2675 555
rect 2833 488 2879 534
rect 3289 515 3335 655
rect 3493 515 3539 655
<< polysilicon >>
rect 144 715 244 760
rect 580 720 3028 760
rect 412 628 512 672
rect 580 628 680 720
rect 748 628 848 672
rect 972 628 1072 672
rect 1196 628 1296 672
rect 1488 628 1588 720
rect 1692 628 1792 672
rect 2100 612 2200 720
rect 144 421 244 472
rect 144 288 185 421
rect 124 280 185 288
rect 231 280 244 421
rect 412 412 512 496
rect 412 366 453 412
rect 499 366 512 412
rect 412 288 512 366
rect 580 288 680 496
rect 748 370 848 496
rect 748 324 789 370
rect 835 324 848 370
rect 748 288 848 324
rect 972 463 1072 496
rect 972 417 1013 463
rect 1059 417 1072 463
rect 972 288 1072 417
rect 1196 288 1296 496
rect 124 232 244 280
rect 392 232 512 288
rect 560 232 680 288
rect 728 232 848 288
rect 952 232 1072 288
rect 1176 232 1296 288
rect 1488 288 1588 496
rect 1692 370 1792 496
rect 2392 612 2492 656
rect 2704 612 2804 656
rect 2928 612 3028 720
rect 3364 715 3464 760
rect 3096 612 3196 656
rect 1692 324 1718 370
rect 1764 324 1792 370
rect 1692 311 1792 324
rect 1712 301 1792 311
rect 1488 232 1608 288
rect 1712 232 1832 301
rect 2100 288 2200 472
rect 2080 232 2200 288
rect 2392 288 2492 472
rect 2704 337 2804 472
rect 2704 291 2717 337
rect 2763 291 2804 337
rect 2704 288 2804 291
rect 2928 415 3028 472
rect 2928 369 2969 415
rect 3015 369 3028 415
rect 2928 288 3028 369
rect 3096 288 3196 472
rect 3364 313 3464 472
rect 2392 232 2512 288
rect 2704 232 2824 288
rect 2928 232 3048 288
rect 3096 232 3216 288
rect 3364 267 3377 313
rect 3423 288 3464 313
rect 3423 267 3484 288
rect 3364 232 3484 267
rect 124 46 244 90
rect 392 64 512 156
rect 560 112 680 156
rect 728 112 848 156
rect 952 112 1072 156
rect 1176 64 1296 156
rect 1488 112 1608 156
rect 1712 112 1832 156
rect 2080 112 2200 156
rect 2392 64 2512 156
rect 2704 112 2824 156
rect 2928 112 3048 156
rect 3096 64 3216 156
rect 392 24 3216 64
rect 3364 24 3484 69
<< polycontact >>
rect 185 280 231 421
rect 453 366 499 412
rect 789 324 835 370
rect 1013 417 1059 463
rect 1718 324 1764 370
rect 2717 291 2763 337
rect 2969 369 3015 415
rect 3377 267 3423 313
<< metal1 >>
rect 0 724 3696 844
rect 273 689 319 724
rect 28 663 115 674
rect 28 523 69 663
rect 273 608 319 643
rect 1358 647 1426 724
rect 1358 601 1369 647
rect 1415 601 1426 647
rect 1821 598 1867 724
rect 2262 647 2330 724
rect 2262 601 2273 647
rect 2319 601 2330 647
rect 3289 655 3335 724
rect 1110 558 1178 569
rect 28 218 115 523
rect 185 512 877 558
rect 923 512 942 558
rect 1110 512 1121 558
rect 1167 555 1178 558
rect 1606 558 1674 569
rect 1606 555 1617 558
rect 1167 512 1617 555
rect 1663 512 1674 558
rect 1821 541 1867 552
rect 185 421 231 512
rect 1110 509 1674 512
rect 2014 509 2025 555
rect 2071 509 2521 555
rect 2567 509 2629 555
rect 2675 509 2686 555
rect 2833 534 2880 553
rect 2879 488 2880 534
rect 3289 496 3335 515
rect 3490 655 3566 674
rect 3490 515 3493 655
rect 3539 515 3566 655
rect 2833 463 2880 488
rect 323 412 694 430
rect 1002 417 1013 463
rect 1059 417 2880 463
rect 1002 416 2880 417
rect 323 366 453 412
rect 499 366 694 412
rect 323 354 694 366
rect 778 324 789 370
rect 835 324 1718 370
rect 1764 337 2782 370
rect 1764 324 2717 337
rect 185 278 231 280
rect 2468 291 2717 324
rect 2763 291 2782 337
rect 185 232 923 278
rect 28 172 49 218
rect 95 172 115 218
rect 877 219 923 232
rect 28 122 115 172
rect 273 163 319 174
rect 877 162 923 173
rect 1101 229 1683 275
rect 1101 219 1147 229
rect 1637 219 1683 229
rect 1101 162 1147 173
rect 273 60 319 117
rect 1358 137 1369 183
rect 1415 137 1426 183
rect 2005 229 2422 275
rect 2468 240 2782 291
rect 1637 162 1683 173
rect 1850 172 1861 218
rect 1907 172 1918 218
rect 1358 60 1426 137
rect 1850 60 1918 172
rect 2005 215 2051 229
rect 2376 183 2422 229
rect 2005 154 2051 169
rect 2262 137 2273 183
rect 2319 137 2330 183
rect 2262 60 2330 137
rect 2376 137 2585 183
rect 2631 137 2642 183
rect 2376 136 2642 137
rect 2708 110 2782 240
rect 2834 313 2880 416
rect 2928 415 3414 430
rect 2928 369 2969 415
rect 3015 369 3414 415
rect 2928 359 3414 369
rect 2834 267 3377 313
rect 3423 267 3440 313
rect 2834 215 2899 267
rect 2834 169 2853 215
rect 2834 150 2899 169
rect 3490 215 3566 515
rect 3490 169 3513 215
rect 3559 169 3566 215
rect 3490 158 3566 169
rect 3289 142 3335 153
rect 3289 60 3335 96
rect 0 -60 3696 60
<< labels >>
flabel metal1 s 2928 359 3414 430 0 FreeSans 600 0 0 0 B
port 2 nsew default input
flabel metal1 s 778 324 2782 370 0 FreeSans 600 0 0 0 CI
port 3 nsew default input
flabel metal1 s 3490 158 3566 674 0 FreeSans 600 0 0 0 CO
port 4 nsew default output
flabel metal1 s 28 122 115 674 0 FreeSans 600 0 0 0 S
port 5 nsew default output
flabel metal1 s 0 724 3696 844 0 FreeSans 600 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1850 183 1918 218 0 FreeSans 600 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 323 354 694 430 0 FreeSans 600 0 0 0 A
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 2468 240 2782 324 1 CI
port 3 nsew default input
rlabel metal1 s 2708 110 2782 240 1 CI
port 3 nsew default input
rlabel metal1 s 3289 608 3335 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2262 608 2330 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1821 608 1867 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1358 608 1426 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 608 319 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3289 601 3335 608 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2262 601 2330 608 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1821 601 1867 608 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1358 601 1426 608 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3289 541 3335 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1821 541 1867 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3289 496 3335 541 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2262 174 2330 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1850 174 1918 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1358 174 1426 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2262 153 2330 174 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1850 153 1918 174 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1358 153 1426 174 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 153 319 174 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3289 60 3335 153 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2262 60 2330 153 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1850 60 1918 153 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1358 60 1426 153 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 153 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3696 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3696 784
string GDS_END 1172912
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1166226
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
