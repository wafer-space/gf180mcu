magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< metal3 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
<< metal4 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
<< metal5 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
use GF_NI_FILLNC_0  GF_NI_FILLNC_0_0
timestamp 1755724134
transform 1 0 0 0 1 0
box -32 13097 52 69968
<< labels >>
rlabel metal3 s 0 63600 20 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 63600 20 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 62000 20 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 20 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 68400 20 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 20 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 20 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 20 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 20 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 20 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 20 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 20 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 20 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 20 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 66800 20 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 20 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 20 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 20 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 20 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 20 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 20 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 20 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 20 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 20 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 20 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 20 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 63600 20 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 49200 20 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 62000 20 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 50800 20 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 65200 20 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 20 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 20 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 20 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 20 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 20 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 20 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 20 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 68400 20 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 65200 20 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 58800 20 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 20 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 20 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 20 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 20 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 20 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 20 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 20 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 20 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 20 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 66800 20 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 58800 20 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 49200 20 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 20 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 50800 20 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 20 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 60400 20 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 57200 20 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 46000 20 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 39600 20 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 25200 20 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 20400 20 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 17200 20 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 14000 20 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 20 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 20 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 55600 20 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 54000 20 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 52400 20 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 42800 20 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 41200 20 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 36400 20 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 33200 20 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 30000 20 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 26800 20 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 23600 20 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 20 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 20 25000 4 DVDD
port 1 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 20 70000
string GDS_END 17631666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17626542
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
