magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 352 758 870
<< pwell >>
rect -86 -86 758 352
<< metal1 >>
rect 0 724 672 844
rect 49 506 95 724
rect 141 236 202 664
rect 477 536 533 676
rect 248 472 533 536
rect 49 60 95 189
rect 248 120 319 472
rect 365 358 571 426
rect 365 120 426 358
rect 497 60 543 218
rect 0 -60 672 60
<< labels >>
rlabel metal1 s 365 120 426 358 6 A1
port 1 nsew default input
rlabel metal1 s 365 358 571 426 6 A1
port 1 nsew default input
rlabel metal1 s 141 236 202 664 6 A2
port 2 nsew default input
rlabel metal1 s 248 120 319 472 6 ZN
port 3 nsew default output
rlabel metal1 s 248 472 533 536 6 ZN
port 3 nsew default output
rlabel metal1 s 477 536 533 676 6 ZN
port 3 nsew default output
rlabel metal1 s 49 506 95 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 724 672 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s -86 352 758 870 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 758 352 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -60 672 60 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 218 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 189 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 740172
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 737482
<< end >>
