magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< psubdiff >>
rect 70 67883 85816 67902
rect 70 67837 89 67883
rect 135 67837 213 67883
rect 259 67837 337 67883
rect 383 67837 461 67883
rect 507 67837 585 67883
rect 631 67837 709 67883
rect 755 67837 833 67883
rect 879 67837 957 67883
rect 1003 67837 1081 67883
rect 1127 67837 1205 67883
rect 1251 67837 1329 67883
rect 1375 67837 1453 67883
rect 1499 67837 1577 67883
rect 1623 67837 1701 67883
rect 1747 67837 1825 67883
rect 1871 67837 1949 67883
rect 1995 67837 2073 67883
rect 2119 67837 2197 67883
rect 2243 67837 2321 67883
rect 2367 67837 2445 67883
rect 2491 67837 2569 67883
rect 2615 67837 2693 67883
rect 2739 67837 2817 67883
rect 2863 67837 2941 67883
rect 2987 67837 3065 67883
rect 3111 67837 3189 67883
rect 3235 67837 3313 67883
rect 3359 67837 3437 67883
rect 3483 67837 3561 67883
rect 3607 67837 3685 67883
rect 3731 67837 3809 67883
rect 3855 67837 3933 67883
rect 3979 67837 4057 67883
rect 4103 67837 4181 67883
rect 4227 67837 4305 67883
rect 4351 67837 4429 67883
rect 4475 67837 4553 67883
rect 4599 67837 4677 67883
rect 4723 67837 4801 67883
rect 4847 67837 4925 67883
rect 4971 67837 5049 67883
rect 5095 67837 5173 67883
rect 5219 67837 5297 67883
rect 5343 67837 5421 67883
rect 5467 67837 5545 67883
rect 5591 67837 5669 67883
rect 5715 67837 5793 67883
rect 5839 67837 5917 67883
rect 5963 67837 6041 67883
rect 6087 67837 6165 67883
rect 6211 67837 6289 67883
rect 6335 67837 6413 67883
rect 6459 67837 6537 67883
rect 6583 67837 6661 67883
rect 6707 67837 6785 67883
rect 6831 67837 6909 67883
rect 6955 67837 7033 67883
rect 7079 67837 7157 67883
rect 7203 67837 7281 67883
rect 7327 67837 7405 67883
rect 7451 67837 7529 67883
rect 7575 67837 7653 67883
rect 7699 67837 7777 67883
rect 7823 67837 7901 67883
rect 7947 67837 8025 67883
rect 8071 67837 8149 67883
rect 8195 67837 8273 67883
rect 8319 67837 8397 67883
rect 8443 67837 8521 67883
rect 8567 67837 8645 67883
rect 8691 67837 8769 67883
rect 8815 67837 8893 67883
rect 8939 67837 9017 67883
rect 9063 67837 9141 67883
rect 9187 67837 9265 67883
rect 9311 67837 9389 67883
rect 9435 67837 9513 67883
rect 9559 67837 9637 67883
rect 9683 67837 9761 67883
rect 9807 67837 9885 67883
rect 9931 67837 10009 67883
rect 10055 67837 10133 67883
rect 10179 67837 10257 67883
rect 10303 67837 10381 67883
rect 10427 67837 10505 67883
rect 10551 67837 10629 67883
rect 10675 67837 10753 67883
rect 10799 67837 10877 67883
rect 10923 67837 11001 67883
rect 11047 67837 11125 67883
rect 11171 67837 11249 67883
rect 11295 67837 11373 67883
rect 11419 67837 11497 67883
rect 11543 67837 11621 67883
rect 11667 67837 11745 67883
rect 11791 67837 11869 67883
rect 11915 67837 11993 67883
rect 12039 67837 12117 67883
rect 12163 67837 12241 67883
rect 12287 67837 12365 67883
rect 12411 67837 12489 67883
rect 12535 67837 12613 67883
rect 12659 67837 12737 67883
rect 12783 67837 12861 67883
rect 12907 67837 12985 67883
rect 13031 67837 13109 67883
rect 13155 67837 13233 67883
rect 13279 67837 13357 67883
rect 13403 67837 13481 67883
rect 13527 67837 13605 67883
rect 13651 67837 13729 67883
rect 13775 67837 13853 67883
rect 13899 67837 13977 67883
rect 14023 67837 14101 67883
rect 14147 67837 14225 67883
rect 14271 67837 14349 67883
rect 14395 67837 14473 67883
rect 14519 67837 14597 67883
rect 14643 67837 14721 67883
rect 14767 67837 14845 67883
rect 14891 67837 14969 67883
rect 15015 67837 15093 67883
rect 15139 67837 15217 67883
rect 15263 67837 15341 67883
rect 15387 67837 15465 67883
rect 15511 67837 15589 67883
rect 15635 67837 15713 67883
rect 15759 67837 15837 67883
rect 15883 67837 15961 67883
rect 16007 67837 16085 67883
rect 16131 67837 16209 67883
rect 16255 67837 16333 67883
rect 16379 67837 16457 67883
rect 16503 67837 16581 67883
rect 16627 67837 16705 67883
rect 16751 67837 16829 67883
rect 16875 67837 16953 67883
rect 16999 67837 17077 67883
rect 17123 67837 17201 67883
rect 17247 67837 17325 67883
rect 17371 67837 17449 67883
rect 17495 67837 17573 67883
rect 17619 67837 17697 67883
rect 17743 67837 17821 67883
rect 17867 67837 17945 67883
rect 17991 67837 18069 67883
rect 18115 67837 18193 67883
rect 18239 67837 18317 67883
rect 18363 67837 18441 67883
rect 18487 67837 18565 67883
rect 18611 67837 18689 67883
rect 18735 67837 18813 67883
rect 18859 67837 18937 67883
rect 18983 67837 19061 67883
rect 19107 67837 19185 67883
rect 19231 67837 19309 67883
rect 19355 67837 19433 67883
rect 19479 67837 19557 67883
rect 19603 67837 19681 67883
rect 19727 67837 19805 67883
rect 19851 67837 19929 67883
rect 19975 67837 20053 67883
rect 20099 67837 20177 67883
rect 20223 67837 20301 67883
rect 20347 67837 20425 67883
rect 20471 67837 20549 67883
rect 20595 67837 20673 67883
rect 20719 67837 20797 67883
rect 20843 67837 20921 67883
rect 20967 67837 21045 67883
rect 21091 67837 21169 67883
rect 21215 67837 21293 67883
rect 21339 67837 21417 67883
rect 21463 67837 21541 67883
rect 21587 67837 21665 67883
rect 21711 67837 21789 67883
rect 21835 67837 21913 67883
rect 21959 67837 22037 67883
rect 22083 67837 22161 67883
rect 22207 67837 22285 67883
rect 22331 67837 22409 67883
rect 22455 67837 22533 67883
rect 22579 67837 22657 67883
rect 22703 67837 22781 67883
rect 22827 67837 22905 67883
rect 22951 67837 23029 67883
rect 23075 67837 23153 67883
rect 23199 67837 23277 67883
rect 23323 67837 23401 67883
rect 23447 67837 23525 67883
rect 23571 67837 23649 67883
rect 23695 67837 23773 67883
rect 23819 67837 23897 67883
rect 23943 67837 24021 67883
rect 24067 67837 24145 67883
rect 24191 67837 24269 67883
rect 24315 67837 24393 67883
rect 24439 67837 24517 67883
rect 24563 67837 24641 67883
rect 24687 67837 24765 67883
rect 24811 67837 24889 67883
rect 24935 67837 25013 67883
rect 25059 67837 25137 67883
rect 25183 67837 25261 67883
rect 25307 67837 25385 67883
rect 25431 67837 25509 67883
rect 25555 67837 25633 67883
rect 25679 67837 25757 67883
rect 25803 67837 25881 67883
rect 25927 67837 26005 67883
rect 26051 67837 26129 67883
rect 26175 67837 26253 67883
rect 26299 67837 26377 67883
rect 26423 67837 26501 67883
rect 26547 67837 26625 67883
rect 26671 67837 26749 67883
rect 26795 67837 26873 67883
rect 26919 67837 26997 67883
rect 27043 67837 27121 67883
rect 27167 67837 27245 67883
rect 27291 67837 27369 67883
rect 27415 67837 27493 67883
rect 27539 67837 27617 67883
rect 27663 67837 27741 67883
rect 27787 67837 27865 67883
rect 27911 67837 27989 67883
rect 28035 67837 28113 67883
rect 28159 67837 28237 67883
rect 28283 67837 28361 67883
rect 28407 67837 28485 67883
rect 28531 67837 28609 67883
rect 28655 67837 28733 67883
rect 28779 67837 28857 67883
rect 28903 67837 28981 67883
rect 29027 67837 29105 67883
rect 29151 67837 29229 67883
rect 29275 67837 29353 67883
rect 29399 67837 29477 67883
rect 29523 67837 29601 67883
rect 29647 67837 29725 67883
rect 29771 67837 29849 67883
rect 29895 67837 29973 67883
rect 30019 67837 30097 67883
rect 30143 67837 30221 67883
rect 30267 67837 30345 67883
rect 30391 67837 30469 67883
rect 30515 67837 30593 67883
rect 30639 67837 30717 67883
rect 30763 67837 30841 67883
rect 30887 67837 30965 67883
rect 31011 67837 31089 67883
rect 31135 67837 31213 67883
rect 31259 67837 31337 67883
rect 31383 67837 31461 67883
rect 31507 67837 31585 67883
rect 31631 67837 31709 67883
rect 31755 67837 31833 67883
rect 31879 67837 31957 67883
rect 32003 67837 32081 67883
rect 32127 67837 32205 67883
rect 32251 67837 32329 67883
rect 32375 67837 32453 67883
rect 32499 67837 32577 67883
rect 32623 67837 32701 67883
rect 32747 67837 32825 67883
rect 32871 67837 32949 67883
rect 32995 67837 33073 67883
rect 33119 67837 33197 67883
rect 33243 67837 33321 67883
rect 33367 67837 33445 67883
rect 33491 67837 33569 67883
rect 33615 67837 33693 67883
rect 33739 67837 33817 67883
rect 33863 67837 33941 67883
rect 33987 67837 34065 67883
rect 34111 67837 34189 67883
rect 34235 67837 34313 67883
rect 34359 67837 34437 67883
rect 34483 67837 34561 67883
rect 34607 67837 34685 67883
rect 34731 67837 34809 67883
rect 34855 67837 34933 67883
rect 34979 67837 35057 67883
rect 35103 67837 35181 67883
rect 35227 67837 35305 67883
rect 35351 67837 35429 67883
rect 35475 67837 35553 67883
rect 35599 67837 35677 67883
rect 35723 67837 35801 67883
rect 35847 67837 35925 67883
rect 35971 67837 36049 67883
rect 36095 67837 36173 67883
rect 36219 67837 36297 67883
rect 36343 67837 36421 67883
rect 36467 67837 36545 67883
rect 36591 67837 36669 67883
rect 36715 67837 36793 67883
rect 36839 67837 36917 67883
rect 36963 67837 37041 67883
rect 37087 67837 37165 67883
rect 37211 67837 37289 67883
rect 37335 67837 37413 67883
rect 37459 67837 37537 67883
rect 37583 67837 37661 67883
rect 37707 67837 37785 67883
rect 37831 67837 37909 67883
rect 37955 67837 38033 67883
rect 38079 67837 38157 67883
rect 38203 67837 38281 67883
rect 38327 67837 38405 67883
rect 38451 67837 38529 67883
rect 38575 67837 38653 67883
rect 38699 67837 38777 67883
rect 38823 67837 38901 67883
rect 38947 67837 39025 67883
rect 39071 67837 39149 67883
rect 39195 67837 39273 67883
rect 39319 67837 39397 67883
rect 39443 67837 39521 67883
rect 39567 67837 39645 67883
rect 39691 67837 39769 67883
rect 39815 67837 39893 67883
rect 39939 67837 40017 67883
rect 40063 67837 40141 67883
rect 40187 67837 40265 67883
rect 40311 67837 40389 67883
rect 40435 67837 40513 67883
rect 40559 67837 40637 67883
rect 40683 67837 40761 67883
rect 40807 67837 40885 67883
rect 40931 67837 41009 67883
rect 41055 67837 41133 67883
rect 41179 67837 41257 67883
rect 41303 67837 41381 67883
rect 41427 67837 41505 67883
rect 41551 67837 41629 67883
rect 41675 67837 41753 67883
rect 41799 67837 41877 67883
rect 41923 67837 42001 67883
rect 42047 67837 42125 67883
rect 42171 67837 42249 67883
rect 42295 67837 42373 67883
rect 42419 67837 42497 67883
rect 42543 67837 42621 67883
rect 42667 67837 42745 67883
rect 42791 67837 42869 67883
rect 42915 67837 42993 67883
rect 43039 67837 43117 67883
rect 43163 67837 43241 67883
rect 43287 67837 43365 67883
rect 43411 67837 43489 67883
rect 43535 67837 43613 67883
rect 43659 67837 43737 67883
rect 43783 67837 43861 67883
rect 43907 67837 43985 67883
rect 44031 67837 44109 67883
rect 44155 67837 44233 67883
rect 44279 67837 44357 67883
rect 44403 67837 44481 67883
rect 44527 67837 44605 67883
rect 44651 67837 44729 67883
rect 44775 67837 44853 67883
rect 44899 67837 44977 67883
rect 45023 67837 45101 67883
rect 45147 67837 45225 67883
rect 45271 67837 45349 67883
rect 45395 67837 45473 67883
rect 45519 67837 45597 67883
rect 45643 67837 45721 67883
rect 45767 67837 45845 67883
rect 45891 67837 45969 67883
rect 46015 67837 46093 67883
rect 46139 67837 46217 67883
rect 46263 67837 46341 67883
rect 46387 67837 46465 67883
rect 46511 67837 46589 67883
rect 46635 67837 46713 67883
rect 46759 67837 46837 67883
rect 46883 67837 46961 67883
rect 47007 67837 47085 67883
rect 47131 67837 47209 67883
rect 47255 67837 47333 67883
rect 47379 67837 47457 67883
rect 47503 67837 47581 67883
rect 47627 67837 47705 67883
rect 47751 67837 47829 67883
rect 47875 67837 47953 67883
rect 47999 67837 48077 67883
rect 48123 67837 48201 67883
rect 48247 67837 48325 67883
rect 48371 67837 48449 67883
rect 48495 67837 48573 67883
rect 48619 67837 48697 67883
rect 48743 67837 48821 67883
rect 48867 67837 48945 67883
rect 48991 67837 49069 67883
rect 49115 67837 49193 67883
rect 49239 67837 49317 67883
rect 49363 67837 49441 67883
rect 49487 67837 49565 67883
rect 49611 67837 49689 67883
rect 49735 67837 49813 67883
rect 49859 67837 49937 67883
rect 49983 67837 50061 67883
rect 50107 67837 50185 67883
rect 50231 67837 50309 67883
rect 50355 67837 50433 67883
rect 50479 67837 50557 67883
rect 50603 67837 50681 67883
rect 50727 67837 50805 67883
rect 50851 67837 50929 67883
rect 50975 67837 51053 67883
rect 51099 67837 51177 67883
rect 51223 67837 51301 67883
rect 51347 67837 51425 67883
rect 51471 67837 51549 67883
rect 51595 67837 51673 67883
rect 51719 67837 51797 67883
rect 51843 67837 51921 67883
rect 51967 67837 52045 67883
rect 52091 67837 52169 67883
rect 52215 67837 52293 67883
rect 52339 67837 52417 67883
rect 52463 67837 52541 67883
rect 52587 67837 52665 67883
rect 52711 67837 52789 67883
rect 52835 67837 52913 67883
rect 52959 67837 53037 67883
rect 53083 67837 53161 67883
rect 53207 67837 53285 67883
rect 53331 67837 53409 67883
rect 53455 67837 53533 67883
rect 53579 67837 53657 67883
rect 53703 67837 53781 67883
rect 53827 67837 53905 67883
rect 53951 67837 54029 67883
rect 54075 67837 54153 67883
rect 54199 67837 54277 67883
rect 54323 67837 54401 67883
rect 54447 67837 54525 67883
rect 54571 67837 54649 67883
rect 54695 67837 54773 67883
rect 54819 67837 54897 67883
rect 54943 67837 55021 67883
rect 55067 67837 55145 67883
rect 55191 67837 55269 67883
rect 55315 67837 55393 67883
rect 55439 67837 55517 67883
rect 55563 67837 55641 67883
rect 55687 67837 55765 67883
rect 55811 67837 55889 67883
rect 55935 67837 56013 67883
rect 56059 67837 56137 67883
rect 56183 67837 56261 67883
rect 56307 67837 56385 67883
rect 56431 67837 56509 67883
rect 56555 67837 56633 67883
rect 56679 67837 56757 67883
rect 56803 67837 56881 67883
rect 56927 67837 57005 67883
rect 57051 67837 57129 67883
rect 57175 67837 57253 67883
rect 57299 67837 57377 67883
rect 57423 67837 57501 67883
rect 57547 67837 57625 67883
rect 57671 67837 57749 67883
rect 57795 67837 57873 67883
rect 57919 67837 57997 67883
rect 58043 67837 58121 67883
rect 58167 67837 58245 67883
rect 58291 67837 58369 67883
rect 58415 67837 58493 67883
rect 58539 67837 58617 67883
rect 58663 67837 58741 67883
rect 58787 67837 58865 67883
rect 58911 67837 58989 67883
rect 59035 67837 59113 67883
rect 59159 67837 59237 67883
rect 59283 67837 59361 67883
rect 59407 67837 59485 67883
rect 59531 67837 59609 67883
rect 59655 67837 59733 67883
rect 59779 67837 59857 67883
rect 59903 67837 59981 67883
rect 60027 67837 60105 67883
rect 60151 67837 60229 67883
rect 60275 67837 60353 67883
rect 60399 67837 60477 67883
rect 60523 67837 60601 67883
rect 60647 67837 60725 67883
rect 60771 67837 60849 67883
rect 60895 67837 60973 67883
rect 61019 67837 61097 67883
rect 61143 67837 61221 67883
rect 61267 67837 61345 67883
rect 61391 67837 61469 67883
rect 61515 67837 61593 67883
rect 61639 67837 61717 67883
rect 61763 67837 61841 67883
rect 61887 67837 61965 67883
rect 62011 67837 62089 67883
rect 62135 67837 62213 67883
rect 62259 67837 62337 67883
rect 62383 67837 62461 67883
rect 62507 67837 62585 67883
rect 62631 67837 62709 67883
rect 62755 67837 62833 67883
rect 62879 67837 62957 67883
rect 63003 67837 63081 67883
rect 63127 67837 63205 67883
rect 63251 67837 63329 67883
rect 63375 67837 63453 67883
rect 63499 67837 63577 67883
rect 63623 67837 63701 67883
rect 63747 67837 63825 67883
rect 63871 67837 63949 67883
rect 63995 67837 64073 67883
rect 64119 67837 64197 67883
rect 64243 67837 64321 67883
rect 64367 67837 64445 67883
rect 64491 67837 64569 67883
rect 64615 67837 64693 67883
rect 64739 67837 64817 67883
rect 64863 67837 64941 67883
rect 64987 67837 65065 67883
rect 65111 67837 65189 67883
rect 65235 67837 65313 67883
rect 65359 67837 65437 67883
rect 65483 67837 65561 67883
rect 65607 67837 65685 67883
rect 65731 67837 65809 67883
rect 65855 67837 65933 67883
rect 65979 67837 66057 67883
rect 66103 67837 66181 67883
rect 66227 67837 66305 67883
rect 66351 67837 66429 67883
rect 66475 67837 66553 67883
rect 66599 67837 66677 67883
rect 66723 67837 66801 67883
rect 66847 67837 66925 67883
rect 66971 67837 67049 67883
rect 67095 67837 67173 67883
rect 67219 67837 67297 67883
rect 67343 67837 67421 67883
rect 67467 67837 67545 67883
rect 67591 67837 67669 67883
rect 67715 67837 67793 67883
rect 67839 67837 67917 67883
rect 67963 67837 68041 67883
rect 68087 67837 68165 67883
rect 68211 67837 68289 67883
rect 68335 67837 68413 67883
rect 68459 67837 68537 67883
rect 68583 67837 68661 67883
rect 68707 67837 68785 67883
rect 68831 67837 68909 67883
rect 68955 67837 69033 67883
rect 69079 67837 69157 67883
rect 69203 67837 69281 67883
rect 69327 67837 69405 67883
rect 69451 67837 69529 67883
rect 69575 67837 69653 67883
rect 69699 67837 69777 67883
rect 69823 67837 69901 67883
rect 69947 67837 70025 67883
rect 70071 67837 70149 67883
rect 70195 67837 70273 67883
rect 70319 67837 70397 67883
rect 70443 67837 70521 67883
rect 70567 67837 70645 67883
rect 70691 67837 70769 67883
rect 70815 67837 70893 67883
rect 70939 67837 71017 67883
rect 71063 67837 71141 67883
rect 71187 67837 71265 67883
rect 71311 67837 71389 67883
rect 71435 67837 71513 67883
rect 71559 67837 71637 67883
rect 71683 67837 71761 67883
rect 71807 67837 71885 67883
rect 71931 67837 72009 67883
rect 72055 67837 72133 67883
rect 72179 67837 72257 67883
rect 72303 67837 72381 67883
rect 72427 67837 72505 67883
rect 72551 67837 72629 67883
rect 72675 67837 72753 67883
rect 72799 67837 72877 67883
rect 72923 67837 73001 67883
rect 73047 67837 73125 67883
rect 73171 67837 73249 67883
rect 73295 67837 73373 67883
rect 73419 67837 73497 67883
rect 73543 67837 73621 67883
rect 73667 67837 73745 67883
rect 73791 67837 73869 67883
rect 73915 67837 73993 67883
rect 74039 67837 74117 67883
rect 74163 67837 74241 67883
rect 74287 67837 74365 67883
rect 74411 67837 74489 67883
rect 74535 67837 74613 67883
rect 74659 67837 74737 67883
rect 74783 67837 74861 67883
rect 74907 67837 74985 67883
rect 75031 67837 75109 67883
rect 75155 67837 75233 67883
rect 75279 67837 75357 67883
rect 75403 67837 75481 67883
rect 75527 67837 75605 67883
rect 75651 67837 75729 67883
rect 75775 67837 75853 67883
rect 75899 67837 75977 67883
rect 76023 67837 76101 67883
rect 76147 67837 76225 67883
rect 76271 67837 76349 67883
rect 76395 67837 76473 67883
rect 76519 67837 76597 67883
rect 76643 67837 76721 67883
rect 76767 67837 76845 67883
rect 76891 67837 76969 67883
rect 77015 67837 77093 67883
rect 77139 67837 77217 67883
rect 77263 67837 77341 67883
rect 77387 67837 77465 67883
rect 77511 67837 77589 67883
rect 77635 67837 77713 67883
rect 77759 67837 77837 67883
rect 77883 67837 77961 67883
rect 78007 67837 78085 67883
rect 78131 67837 78209 67883
rect 78255 67837 78333 67883
rect 78379 67837 78457 67883
rect 78503 67837 78581 67883
rect 78627 67837 78705 67883
rect 78751 67837 78829 67883
rect 78875 67837 78953 67883
rect 78999 67837 79077 67883
rect 79123 67837 79201 67883
rect 79247 67837 79325 67883
rect 79371 67837 79449 67883
rect 79495 67837 79573 67883
rect 79619 67837 79697 67883
rect 79743 67837 79821 67883
rect 79867 67837 79945 67883
rect 79991 67837 80069 67883
rect 80115 67837 80193 67883
rect 80239 67837 80317 67883
rect 80363 67837 80441 67883
rect 80487 67837 80565 67883
rect 80611 67837 80689 67883
rect 80735 67837 80813 67883
rect 80859 67837 80937 67883
rect 80983 67837 81061 67883
rect 81107 67837 81185 67883
rect 81231 67837 81309 67883
rect 81355 67837 81433 67883
rect 81479 67837 81557 67883
rect 81603 67837 81681 67883
rect 81727 67837 81805 67883
rect 81851 67837 81929 67883
rect 81975 67837 82053 67883
rect 82099 67837 82177 67883
rect 82223 67837 82301 67883
rect 82347 67837 82425 67883
rect 82471 67837 82549 67883
rect 82595 67837 82673 67883
rect 82719 67837 82797 67883
rect 82843 67837 82921 67883
rect 82967 67837 83045 67883
rect 83091 67837 83169 67883
rect 83215 67837 83293 67883
rect 83339 67837 83417 67883
rect 83463 67837 83541 67883
rect 83587 67837 83665 67883
rect 83711 67837 83789 67883
rect 83835 67837 83913 67883
rect 83959 67837 84037 67883
rect 84083 67837 84161 67883
rect 84207 67837 84285 67883
rect 84331 67837 84409 67883
rect 84455 67837 84533 67883
rect 84579 67837 84657 67883
rect 84703 67837 84781 67883
rect 84827 67837 84905 67883
rect 84951 67837 85029 67883
rect 85075 67837 85153 67883
rect 85199 67837 85277 67883
rect 85323 67837 85401 67883
rect 85447 67837 85525 67883
rect 85571 67837 85649 67883
rect 85695 67837 85816 67883
rect 70 67759 85816 67837
rect 70 67713 89 67759
rect 135 67713 213 67759
rect 259 67713 337 67759
rect 383 67713 461 67759
rect 507 67713 585 67759
rect 631 67713 709 67759
rect 755 67713 833 67759
rect 879 67713 957 67759
rect 1003 67713 1081 67759
rect 1127 67713 1205 67759
rect 1251 67713 1329 67759
rect 1375 67713 1453 67759
rect 1499 67713 1577 67759
rect 1623 67713 1701 67759
rect 1747 67713 1825 67759
rect 1871 67713 1949 67759
rect 1995 67713 2073 67759
rect 2119 67713 2197 67759
rect 2243 67713 2321 67759
rect 2367 67713 2445 67759
rect 2491 67713 2569 67759
rect 2615 67713 2693 67759
rect 2739 67713 2817 67759
rect 2863 67713 2941 67759
rect 2987 67713 3065 67759
rect 3111 67713 3189 67759
rect 3235 67713 3313 67759
rect 3359 67713 3437 67759
rect 3483 67713 3561 67759
rect 3607 67713 3685 67759
rect 3731 67713 3809 67759
rect 3855 67713 3933 67759
rect 3979 67713 4057 67759
rect 4103 67713 4181 67759
rect 4227 67713 4305 67759
rect 4351 67713 4429 67759
rect 4475 67713 4553 67759
rect 4599 67713 4677 67759
rect 4723 67713 4801 67759
rect 4847 67713 4925 67759
rect 4971 67713 5049 67759
rect 5095 67713 5173 67759
rect 5219 67713 5297 67759
rect 5343 67713 5421 67759
rect 5467 67713 5545 67759
rect 5591 67713 5669 67759
rect 5715 67713 5793 67759
rect 5839 67713 5917 67759
rect 5963 67713 6041 67759
rect 6087 67713 6165 67759
rect 6211 67713 6289 67759
rect 6335 67713 6413 67759
rect 6459 67713 6537 67759
rect 6583 67713 6661 67759
rect 6707 67713 6785 67759
rect 6831 67713 6909 67759
rect 6955 67713 7033 67759
rect 7079 67713 7157 67759
rect 7203 67713 7281 67759
rect 7327 67713 7405 67759
rect 7451 67713 7529 67759
rect 7575 67713 7653 67759
rect 7699 67713 7777 67759
rect 7823 67713 7901 67759
rect 7947 67713 8025 67759
rect 8071 67713 8149 67759
rect 8195 67713 8273 67759
rect 8319 67713 8397 67759
rect 8443 67713 8521 67759
rect 8567 67713 8645 67759
rect 8691 67713 8769 67759
rect 8815 67713 8893 67759
rect 8939 67713 9017 67759
rect 9063 67713 9141 67759
rect 9187 67713 9265 67759
rect 9311 67713 9389 67759
rect 9435 67713 9513 67759
rect 9559 67713 9637 67759
rect 9683 67713 9761 67759
rect 9807 67713 9885 67759
rect 9931 67713 10009 67759
rect 10055 67713 10133 67759
rect 10179 67713 10257 67759
rect 10303 67713 10381 67759
rect 10427 67713 10505 67759
rect 10551 67713 10629 67759
rect 10675 67713 10753 67759
rect 10799 67713 10877 67759
rect 10923 67713 11001 67759
rect 11047 67713 11125 67759
rect 11171 67713 11249 67759
rect 11295 67713 11373 67759
rect 11419 67713 11497 67759
rect 11543 67713 11621 67759
rect 11667 67713 11745 67759
rect 11791 67713 11869 67759
rect 11915 67713 11993 67759
rect 12039 67713 12117 67759
rect 12163 67713 12241 67759
rect 12287 67713 12365 67759
rect 12411 67713 12489 67759
rect 12535 67713 12613 67759
rect 12659 67713 12737 67759
rect 12783 67713 12861 67759
rect 12907 67713 12985 67759
rect 13031 67713 13109 67759
rect 13155 67713 13233 67759
rect 13279 67713 13357 67759
rect 13403 67713 13481 67759
rect 13527 67713 13605 67759
rect 13651 67713 13729 67759
rect 13775 67713 13853 67759
rect 13899 67713 13977 67759
rect 14023 67713 14101 67759
rect 14147 67713 14225 67759
rect 14271 67713 14349 67759
rect 14395 67713 14473 67759
rect 14519 67713 14597 67759
rect 14643 67713 14721 67759
rect 14767 67713 14845 67759
rect 14891 67713 14969 67759
rect 15015 67713 15093 67759
rect 15139 67713 15217 67759
rect 15263 67713 15341 67759
rect 15387 67713 15465 67759
rect 15511 67713 15589 67759
rect 15635 67713 15713 67759
rect 15759 67713 15837 67759
rect 15883 67713 15961 67759
rect 16007 67713 16085 67759
rect 16131 67713 16209 67759
rect 16255 67713 16333 67759
rect 16379 67713 16457 67759
rect 16503 67713 16581 67759
rect 16627 67713 16705 67759
rect 16751 67713 16829 67759
rect 16875 67713 16953 67759
rect 16999 67713 17077 67759
rect 17123 67713 17201 67759
rect 17247 67713 17325 67759
rect 17371 67713 17449 67759
rect 17495 67713 17573 67759
rect 17619 67713 17697 67759
rect 17743 67713 17821 67759
rect 17867 67713 17945 67759
rect 17991 67713 18069 67759
rect 18115 67713 18193 67759
rect 18239 67713 18317 67759
rect 18363 67713 18441 67759
rect 18487 67713 18565 67759
rect 18611 67713 18689 67759
rect 18735 67713 18813 67759
rect 18859 67713 18937 67759
rect 18983 67713 19061 67759
rect 19107 67713 19185 67759
rect 19231 67713 19309 67759
rect 19355 67713 19433 67759
rect 19479 67713 19557 67759
rect 19603 67713 19681 67759
rect 19727 67713 19805 67759
rect 19851 67713 19929 67759
rect 19975 67713 20053 67759
rect 20099 67713 20177 67759
rect 20223 67713 20301 67759
rect 20347 67713 20425 67759
rect 20471 67713 20549 67759
rect 20595 67713 20673 67759
rect 20719 67713 20797 67759
rect 20843 67713 20921 67759
rect 20967 67713 21045 67759
rect 21091 67713 21169 67759
rect 21215 67713 21293 67759
rect 21339 67713 21417 67759
rect 21463 67713 21541 67759
rect 21587 67713 21665 67759
rect 21711 67713 21789 67759
rect 21835 67713 21913 67759
rect 21959 67713 22037 67759
rect 22083 67713 22161 67759
rect 22207 67713 22285 67759
rect 22331 67713 22409 67759
rect 22455 67713 22533 67759
rect 22579 67713 22657 67759
rect 22703 67713 22781 67759
rect 22827 67713 22905 67759
rect 22951 67713 23029 67759
rect 23075 67713 23153 67759
rect 23199 67713 23277 67759
rect 23323 67713 23401 67759
rect 23447 67713 23525 67759
rect 23571 67713 23649 67759
rect 23695 67713 23773 67759
rect 23819 67713 23897 67759
rect 23943 67713 24021 67759
rect 24067 67713 24145 67759
rect 24191 67713 24269 67759
rect 24315 67713 24393 67759
rect 24439 67713 24517 67759
rect 24563 67713 24641 67759
rect 24687 67713 24765 67759
rect 24811 67713 24889 67759
rect 24935 67713 25013 67759
rect 25059 67713 25137 67759
rect 25183 67713 25261 67759
rect 25307 67713 25385 67759
rect 25431 67713 25509 67759
rect 25555 67713 25633 67759
rect 25679 67713 25757 67759
rect 25803 67713 25881 67759
rect 25927 67713 26005 67759
rect 26051 67713 26129 67759
rect 26175 67713 26253 67759
rect 26299 67713 26377 67759
rect 26423 67713 26501 67759
rect 26547 67713 26625 67759
rect 26671 67713 26749 67759
rect 26795 67713 26873 67759
rect 26919 67713 26997 67759
rect 27043 67713 27121 67759
rect 27167 67713 27245 67759
rect 27291 67713 27369 67759
rect 27415 67713 27493 67759
rect 27539 67713 27617 67759
rect 27663 67713 27741 67759
rect 27787 67713 27865 67759
rect 27911 67713 27989 67759
rect 28035 67713 28113 67759
rect 28159 67713 28237 67759
rect 28283 67713 28361 67759
rect 28407 67713 28485 67759
rect 28531 67713 28609 67759
rect 28655 67713 28733 67759
rect 28779 67713 28857 67759
rect 28903 67713 28981 67759
rect 29027 67713 29105 67759
rect 29151 67713 29229 67759
rect 29275 67713 29353 67759
rect 29399 67713 29477 67759
rect 29523 67713 29601 67759
rect 29647 67713 29725 67759
rect 29771 67713 29849 67759
rect 29895 67713 29973 67759
rect 30019 67713 30097 67759
rect 30143 67713 30221 67759
rect 30267 67713 30345 67759
rect 30391 67713 30469 67759
rect 30515 67713 30593 67759
rect 30639 67713 30717 67759
rect 30763 67713 30841 67759
rect 30887 67713 30965 67759
rect 31011 67713 31089 67759
rect 31135 67713 31213 67759
rect 31259 67713 31337 67759
rect 31383 67713 31461 67759
rect 31507 67713 31585 67759
rect 31631 67713 31709 67759
rect 31755 67713 31833 67759
rect 31879 67713 31957 67759
rect 32003 67713 32081 67759
rect 32127 67713 32205 67759
rect 32251 67713 32329 67759
rect 32375 67713 32453 67759
rect 32499 67713 32577 67759
rect 32623 67713 32701 67759
rect 32747 67713 32825 67759
rect 32871 67713 32949 67759
rect 32995 67713 33073 67759
rect 33119 67713 33197 67759
rect 33243 67713 33321 67759
rect 33367 67713 33445 67759
rect 33491 67713 33569 67759
rect 33615 67713 33693 67759
rect 33739 67713 33817 67759
rect 33863 67713 33941 67759
rect 33987 67713 34065 67759
rect 34111 67713 34189 67759
rect 34235 67713 34313 67759
rect 34359 67713 34437 67759
rect 34483 67713 34561 67759
rect 34607 67713 34685 67759
rect 34731 67713 34809 67759
rect 34855 67713 34933 67759
rect 34979 67713 35057 67759
rect 35103 67713 35181 67759
rect 35227 67713 35305 67759
rect 35351 67713 35429 67759
rect 35475 67713 35553 67759
rect 35599 67713 35677 67759
rect 35723 67713 35801 67759
rect 35847 67713 35925 67759
rect 35971 67713 36049 67759
rect 36095 67713 36173 67759
rect 36219 67713 36297 67759
rect 36343 67713 36421 67759
rect 36467 67713 36545 67759
rect 36591 67713 36669 67759
rect 36715 67713 36793 67759
rect 36839 67713 36917 67759
rect 36963 67713 37041 67759
rect 37087 67713 37165 67759
rect 37211 67713 37289 67759
rect 37335 67713 37413 67759
rect 37459 67713 37537 67759
rect 37583 67713 37661 67759
rect 37707 67713 37785 67759
rect 37831 67713 37909 67759
rect 37955 67713 38033 67759
rect 38079 67713 38157 67759
rect 38203 67713 38281 67759
rect 38327 67713 38405 67759
rect 38451 67713 38529 67759
rect 38575 67713 38653 67759
rect 38699 67713 38777 67759
rect 38823 67713 38901 67759
rect 38947 67713 39025 67759
rect 39071 67713 39149 67759
rect 39195 67713 39273 67759
rect 39319 67713 39397 67759
rect 39443 67713 39521 67759
rect 39567 67713 39645 67759
rect 39691 67713 39769 67759
rect 39815 67713 39893 67759
rect 39939 67713 40017 67759
rect 40063 67713 40141 67759
rect 40187 67713 40265 67759
rect 40311 67713 40389 67759
rect 40435 67713 40513 67759
rect 40559 67713 40637 67759
rect 40683 67713 40761 67759
rect 40807 67713 40885 67759
rect 40931 67713 41009 67759
rect 41055 67713 41133 67759
rect 41179 67713 41257 67759
rect 41303 67713 41381 67759
rect 41427 67713 41505 67759
rect 41551 67713 41629 67759
rect 41675 67713 41753 67759
rect 41799 67713 41877 67759
rect 41923 67713 42001 67759
rect 42047 67713 42125 67759
rect 42171 67713 42249 67759
rect 42295 67713 42373 67759
rect 42419 67713 42497 67759
rect 42543 67713 42621 67759
rect 42667 67713 42745 67759
rect 42791 67713 42869 67759
rect 42915 67713 42993 67759
rect 43039 67713 43117 67759
rect 43163 67713 43241 67759
rect 43287 67713 43365 67759
rect 43411 67713 43489 67759
rect 43535 67713 43613 67759
rect 43659 67713 43737 67759
rect 43783 67713 43861 67759
rect 43907 67713 43985 67759
rect 44031 67713 44109 67759
rect 44155 67713 44233 67759
rect 44279 67713 44357 67759
rect 44403 67713 44481 67759
rect 44527 67713 44605 67759
rect 44651 67713 44729 67759
rect 44775 67713 44853 67759
rect 44899 67713 44977 67759
rect 45023 67713 45101 67759
rect 45147 67713 45225 67759
rect 45271 67713 45349 67759
rect 45395 67713 45473 67759
rect 45519 67713 45597 67759
rect 45643 67713 45721 67759
rect 45767 67713 45845 67759
rect 45891 67713 45969 67759
rect 46015 67713 46093 67759
rect 46139 67713 46217 67759
rect 46263 67713 46341 67759
rect 46387 67713 46465 67759
rect 46511 67713 46589 67759
rect 46635 67713 46713 67759
rect 46759 67713 46837 67759
rect 46883 67713 46961 67759
rect 47007 67713 47085 67759
rect 47131 67713 47209 67759
rect 47255 67713 47333 67759
rect 47379 67713 47457 67759
rect 47503 67713 47581 67759
rect 47627 67713 47705 67759
rect 47751 67713 47829 67759
rect 47875 67713 47953 67759
rect 47999 67713 48077 67759
rect 48123 67713 48201 67759
rect 48247 67713 48325 67759
rect 48371 67713 48449 67759
rect 48495 67713 48573 67759
rect 48619 67713 48697 67759
rect 48743 67713 48821 67759
rect 48867 67713 48945 67759
rect 48991 67713 49069 67759
rect 49115 67713 49193 67759
rect 49239 67713 49317 67759
rect 49363 67713 49441 67759
rect 49487 67713 49565 67759
rect 49611 67713 49689 67759
rect 49735 67713 49813 67759
rect 49859 67713 49937 67759
rect 49983 67713 50061 67759
rect 50107 67713 50185 67759
rect 50231 67713 50309 67759
rect 50355 67713 50433 67759
rect 50479 67713 50557 67759
rect 50603 67713 50681 67759
rect 50727 67713 50805 67759
rect 50851 67713 50929 67759
rect 50975 67713 51053 67759
rect 51099 67713 51177 67759
rect 51223 67713 51301 67759
rect 51347 67713 51425 67759
rect 51471 67713 51549 67759
rect 51595 67713 51673 67759
rect 51719 67713 51797 67759
rect 51843 67713 51921 67759
rect 51967 67713 52045 67759
rect 52091 67713 52169 67759
rect 52215 67713 52293 67759
rect 52339 67713 52417 67759
rect 52463 67713 52541 67759
rect 52587 67713 52665 67759
rect 52711 67713 52789 67759
rect 52835 67713 52913 67759
rect 52959 67713 53037 67759
rect 53083 67713 53161 67759
rect 53207 67713 53285 67759
rect 53331 67713 53409 67759
rect 53455 67713 53533 67759
rect 53579 67713 53657 67759
rect 53703 67713 53781 67759
rect 53827 67713 53905 67759
rect 53951 67713 54029 67759
rect 54075 67713 54153 67759
rect 54199 67713 54277 67759
rect 54323 67713 54401 67759
rect 54447 67713 54525 67759
rect 54571 67713 54649 67759
rect 54695 67713 54773 67759
rect 54819 67713 54897 67759
rect 54943 67713 55021 67759
rect 55067 67713 55145 67759
rect 55191 67713 55269 67759
rect 55315 67713 55393 67759
rect 55439 67713 55517 67759
rect 55563 67713 55641 67759
rect 55687 67713 55765 67759
rect 55811 67713 55889 67759
rect 55935 67713 56013 67759
rect 56059 67713 56137 67759
rect 56183 67713 56261 67759
rect 56307 67713 56385 67759
rect 56431 67713 56509 67759
rect 56555 67713 56633 67759
rect 56679 67713 56757 67759
rect 56803 67713 56881 67759
rect 56927 67713 57005 67759
rect 57051 67713 57129 67759
rect 57175 67713 57253 67759
rect 57299 67713 57377 67759
rect 57423 67713 57501 67759
rect 57547 67713 57625 67759
rect 57671 67713 57749 67759
rect 57795 67713 57873 67759
rect 57919 67713 57997 67759
rect 58043 67713 58121 67759
rect 58167 67713 58245 67759
rect 58291 67713 58369 67759
rect 58415 67713 58493 67759
rect 58539 67713 58617 67759
rect 58663 67713 58741 67759
rect 58787 67713 58865 67759
rect 58911 67713 58989 67759
rect 59035 67713 59113 67759
rect 59159 67713 59237 67759
rect 59283 67713 59361 67759
rect 59407 67713 59485 67759
rect 59531 67713 59609 67759
rect 59655 67713 59733 67759
rect 59779 67713 59857 67759
rect 59903 67713 59981 67759
rect 60027 67713 60105 67759
rect 60151 67713 60229 67759
rect 60275 67713 60353 67759
rect 60399 67713 60477 67759
rect 60523 67713 60601 67759
rect 60647 67713 60725 67759
rect 60771 67713 60849 67759
rect 60895 67713 60973 67759
rect 61019 67713 61097 67759
rect 61143 67713 61221 67759
rect 61267 67713 61345 67759
rect 61391 67713 61469 67759
rect 61515 67713 61593 67759
rect 61639 67713 61717 67759
rect 61763 67713 61841 67759
rect 61887 67713 61965 67759
rect 62011 67713 62089 67759
rect 62135 67713 62213 67759
rect 62259 67713 62337 67759
rect 62383 67713 62461 67759
rect 62507 67713 62585 67759
rect 62631 67713 62709 67759
rect 62755 67713 62833 67759
rect 62879 67713 62957 67759
rect 63003 67713 63081 67759
rect 63127 67713 63205 67759
rect 63251 67713 63329 67759
rect 63375 67713 63453 67759
rect 63499 67713 63577 67759
rect 63623 67713 63701 67759
rect 63747 67713 63825 67759
rect 63871 67713 63949 67759
rect 63995 67713 64073 67759
rect 64119 67713 64197 67759
rect 64243 67713 64321 67759
rect 64367 67713 64445 67759
rect 64491 67713 64569 67759
rect 64615 67713 64693 67759
rect 64739 67713 64817 67759
rect 64863 67713 64941 67759
rect 64987 67713 65065 67759
rect 65111 67713 65189 67759
rect 65235 67713 65313 67759
rect 65359 67713 65437 67759
rect 65483 67713 65561 67759
rect 65607 67713 65685 67759
rect 65731 67713 65809 67759
rect 65855 67713 65933 67759
rect 65979 67713 66057 67759
rect 66103 67713 66181 67759
rect 66227 67713 66305 67759
rect 66351 67713 66429 67759
rect 66475 67713 66553 67759
rect 66599 67713 66677 67759
rect 66723 67713 66801 67759
rect 66847 67713 66925 67759
rect 66971 67713 67049 67759
rect 67095 67713 67173 67759
rect 67219 67713 67297 67759
rect 67343 67713 67421 67759
rect 67467 67713 67545 67759
rect 67591 67713 67669 67759
rect 67715 67713 67793 67759
rect 67839 67713 67917 67759
rect 67963 67713 68041 67759
rect 68087 67713 68165 67759
rect 68211 67713 68289 67759
rect 68335 67713 68413 67759
rect 68459 67713 68537 67759
rect 68583 67713 68661 67759
rect 68707 67713 68785 67759
rect 68831 67713 68909 67759
rect 68955 67713 69033 67759
rect 69079 67713 69157 67759
rect 69203 67713 69281 67759
rect 69327 67713 69405 67759
rect 69451 67713 69529 67759
rect 69575 67713 69653 67759
rect 69699 67713 69777 67759
rect 69823 67713 69901 67759
rect 69947 67713 70025 67759
rect 70071 67713 70149 67759
rect 70195 67713 70273 67759
rect 70319 67713 70397 67759
rect 70443 67713 70521 67759
rect 70567 67713 70645 67759
rect 70691 67713 70769 67759
rect 70815 67713 70893 67759
rect 70939 67713 71017 67759
rect 71063 67713 71141 67759
rect 71187 67713 71265 67759
rect 71311 67713 71389 67759
rect 71435 67713 71513 67759
rect 71559 67713 71637 67759
rect 71683 67713 71761 67759
rect 71807 67713 71885 67759
rect 71931 67713 72009 67759
rect 72055 67713 72133 67759
rect 72179 67713 72257 67759
rect 72303 67713 72381 67759
rect 72427 67713 72505 67759
rect 72551 67713 72629 67759
rect 72675 67713 72753 67759
rect 72799 67713 72877 67759
rect 72923 67713 73001 67759
rect 73047 67713 73125 67759
rect 73171 67713 73249 67759
rect 73295 67713 73373 67759
rect 73419 67713 73497 67759
rect 73543 67713 73621 67759
rect 73667 67713 73745 67759
rect 73791 67713 73869 67759
rect 73915 67713 73993 67759
rect 74039 67713 74117 67759
rect 74163 67713 74241 67759
rect 74287 67713 74365 67759
rect 74411 67713 74489 67759
rect 74535 67713 74613 67759
rect 74659 67713 74737 67759
rect 74783 67713 74861 67759
rect 74907 67713 74985 67759
rect 75031 67713 75109 67759
rect 75155 67713 75233 67759
rect 75279 67713 75357 67759
rect 75403 67713 75481 67759
rect 75527 67713 75605 67759
rect 75651 67713 75729 67759
rect 75775 67713 75853 67759
rect 75899 67713 75977 67759
rect 76023 67713 76101 67759
rect 76147 67713 76225 67759
rect 76271 67713 76349 67759
rect 76395 67713 76473 67759
rect 76519 67713 76597 67759
rect 76643 67713 76721 67759
rect 76767 67713 76845 67759
rect 76891 67713 76969 67759
rect 77015 67713 77093 67759
rect 77139 67713 77217 67759
rect 77263 67713 77341 67759
rect 77387 67713 77465 67759
rect 77511 67713 77589 67759
rect 77635 67713 77713 67759
rect 77759 67713 77837 67759
rect 77883 67713 77961 67759
rect 78007 67713 78085 67759
rect 78131 67713 78209 67759
rect 78255 67713 78333 67759
rect 78379 67713 78457 67759
rect 78503 67713 78581 67759
rect 78627 67713 78705 67759
rect 78751 67713 78829 67759
rect 78875 67713 78953 67759
rect 78999 67713 79077 67759
rect 79123 67713 79201 67759
rect 79247 67713 79325 67759
rect 79371 67713 79449 67759
rect 79495 67713 79573 67759
rect 79619 67713 79697 67759
rect 79743 67713 79821 67759
rect 79867 67713 79945 67759
rect 79991 67713 80069 67759
rect 80115 67713 80193 67759
rect 80239 67713 80317 67759
rect 80363 67713 80441 67759
rect 80487 67713 80565 67759
rect 80611 67713 80689 67759
rect 80735 67713 80813 67759
rect 80859 67713 80937 67759
rect 80983 67713 81061 67759
rect 81107 67713 81185 67759
rect 81231 67713 81309 67759
rect 81355 67713 81433 67759
rect 81479 67713 81557 67759
rect 81603 67713 81681 67759
rect 81727 67713 81805 67759
rect 81851 67713 81929 67759
rect 81975 67713 82053 67759
rect 82099 67713 82177 67759
rect 82223 67713 82301 67759
rect 82347 67713 82425 67759
rect 82471 67713 82549 67759
rect 82595 67713 82673 67759
rect 82719 67713 82797 67759
rect 82843 67713 82921 67759
rect 82967 67713 83045 67759
rect 83091 67713 83169 67759
rect 83215 67713 83293 67759
rect 83339 67713 83417 67759
rect 83463 67713 83541 67759
rect 83587 67713 83665 67759
rect 83711 67713 83789 67759
rect 83835 67713 83913 67759
rect 83959 67713 84037 67759
rect 84083 67713 84161 67759
rect 84207 67713 84285 67759
rect 84331 67713 84409 67759
rect 84455 67713 84533 67759
rect 84579 67713 84657 67759
rect 84703 67713 84781 67759
rect 84827 67713 84905 67759
rect 84951 67713 85029 67759
rect 85075 67713 85153 67759
rect 85199 67713 85277 67759
rect 85323 67713 85401 67759
rect 85447 67713 85525 67759
rect 85571 67713 85649 67759
rect 85695 67713 85816 67759
rect 70 67635 85816 67713
rect 70 67589 89 67635
rect 135 67589 213 67635
rect 259 67589 337 67635
rect 383 67589 461 67635
rect 507 67589 585 67635
rect 631 67589 709 67635
rect 755 67589 833 67635
rect 879 67589 957 67635
rect 1003 67589 1081 67635
rect 1127 67589 1205 67635
rect 1251 67589 1329 67635
rect 1375 67589 1453 67635
rect 1499 67589 1577 67635
rect 1623 67589 1701 67635
rect 1747 67589 1825 67635
rect 1871 67589 1949 67635
rect 1995 67589 2073 67635
rect 2119 67589 2197 67635
rect 2243 67589 2321 67635
rect 2367 67589 2445 67635
rect 2491 67589 2569 67635
rect 2615 67589 2693 67635
rect 2739 67589 2817 67635
rect 2863 67589 2941 67635
rect 2987 67589 3065 67635
rect 3111 67589 3189 67635
rect 3235 67589 3313 67635
rect 3359 67589 3437 67635
rect 3483 67589 3561 67635
rect 3607 67589 3685 67635
rect 3731 67589 3809 67635
rect 3855 67589 3933 67635
rect 3979 67589 4057 67635
rect 4103 67589 4181 67635
rect 4227 67589 4305 67635
rect 4351 67589 4429 67635
rect 4475 67589 4553 67635
rect 4599 67589 4677 67635
rect 4723 67589 4801 67635
rect 4847 67589 4925 67635
rect 4971 67589 5049 67635
rect 5095 67589 5173 67635
rect 5219 67589 5297 67635
rect 5343 67589 5421 67635
rect 5467 67589 5545 67635
rect 5591 67589 5669 67635
rect 5715 67589 5793 67635
rect 5839 67589 5917 67635
rect 5963 67589 6041 67635
rect 6087 67589 6165 67635
rect 6211 67589 6289 67635
rect 6335 67589 6413 67635
rect 6459 67589 6537 67635
rect 6583 67589 6661 67635
rect 6707 67589 6785 67635
rect 6831 67589 6909 67635
rect 6955 67589 7033 67635
rect 7079 67589 7157 67635
rect 7203 67589 7281 67635
rect 7327 67589 7405 67635
rect 7451 67589 7529 67635
rect 7575 67589 7653 67635
rect 7699 67589 7777 67635
rect 7823 67589 7901 67635
rect 7947 67589 8025 67635
rect 8071 67589 8149 67635
rect 8195 67589 8273 67635
rect 8319 67589 8397 67635
rect 8443 67589 8521 67635
rect 8567 67589 8645 67635
rect 8691 67589 8769 67635
rect 8815 67589 8893 67635
rect 8939 67589 9017 67635
rect 9063 67589 9141 67635
rect 9187 67589 9265 67635
rect 9311 67589 9389 67635
rect 9435 67589 9513 67635
rect 9559 67589 9637 67635
rect 9683 67589 9761 67635
rect 9807 67589 9885 67635
rect 9931 67589 10009 67635
rect 10055 67589 10133 67635
rect 10179 67589 10257 67635
rect 10303 67589 10381 67635
rect 10427 67589 10505 67635
rect 10551 67589 10629 67635
rect 10675 67589 10753 67635
rect 10799 67589 10877 67635
rect 10923 67589 11001 67635
rect 11047 67589 11125 67635
rect 11171 67589 11249 67635
rect 11295 67589 11373 67635
rect 11419 67589 11497 67635
rect 11543 67589 11621 67635
rect 11667 67589 11745 67635
rect 11791 67589 11869 67635
rect 11915 67589 11993 67635
rect 12039 67589 12117 67635
rect 12163 67589 12241 67635
rect 12287 67589 12365 67635
rect 12411 67589 12489 67635
rect 12535 67589 12613 67635
rect 12659 67589 12737 67635
rect 12783 67589 12861 67635
rect 12907 67589 12985 67635
rect 13031 67589 13109 67635
rect 13155 67589 13233 67635
rect 13279 67589 13357 67635
rect 13403 67589 13481 67635
rect 13527 67589 13605 67635
rect 13651 67589 13729 67635
rect 13775 67589 13853 67635
rect 13899 67589 13977 67635
rect 14023 67589 14101 67635
rect 14147 67589 14225 67635
rect 14271 67589 14349 67635
rect 14395 67589 14473 67635
rect 14519 67589 14597 67635
rect 14643 67589 14721 67635
rect 14767 67589 14845 67635
rect 14891 67589 14969 67635
rect 15015 67589 15093 67635
rect 15139 67589 15217 67635
rect 15263 67589 15341 67635
rect 15387 67589 15465 67635
rect 15511 67589 15589 67635
rect 15635 67589 15713 67635
rect 15759 67589 15837 67635
rect 15883 67589 15961 67635
rect 16007 67589 16085 67635
rect 16131 67589 16209 67635
rect 16255 67589 16333 67635
rect 16379 67589 16457 67635
rect 16503 67589 16581 67635
rect 16627 67589 16705 67635
rect 16751 67589 16829 67635
rect 16875 67589 16953 67635
rect 16999 67589 17077 67635
rect 17123 67589 17201 67635
rect 17247 67589 17325 67635
rect 17371 67589 17449 67635
rect 17495 67589 17573 67635
rect 17619 67589 17697 67635
rect 17743 67589 17821 67635
rect 17867 67589 17945 67635
rect 17991 67589 18069 67635
rect 18115 67589 18193 67635
rect 18239 67589 18317 67635
rect 18363 67589 18441 67635
rect 18487 67589 18565 67635
rect 18611 67589 18689 67635
rect 18735 67589 18813 67635
rect 18859 67589 18937 67635
rect 18983 67589 19061 67635
rect 19107 67589 19185 67635
rect 19231 67589 19309 67635
rect 19355 67589 19433 67635
rect 19479 67589 19557 67635
rect 19603 67589 19681 67635
rect 19727 67589 19805 67635
rect 19851 67589 19929 67635
rect 19975 67589 20053 67635
rect 20099 67589 20177 67635
rect 20223 67589 20301 67635
rect 20347 67589 20425 67635
rect 20471 67589 20549 67635
rect 20595 67589 20673 67635
rect 20719 67589 20797 67635
rect 20843 67589 20921 67635
rect 20967 67589 21045 67635
rect 21091 67589 21169 67635
rect 21215 67589 21293 67635
rect 21339 67589 21417 67635
rect 21463 67589 21541 67635
rect 21587 67589 21665 67635
rect 21711 67589 21789 67635
rect 21835 67589 21913 67635
rect 21959 67589 22037 67635
rect 22083 67589 22161 67635
rect 22207 67589 22285 67635
rect 22331 67589 22409 67635
rect 22455 67589 22533 67635
rect 22579 67589 22657 67635
rect 22703 67589 22781 67635
rect 22827 67589 22905 67635
rect 22951 67589 23029 67635
rect 23075 67589 23153 67635
rect 23199 67589 23277 67635
rect 23323 67589 23401 67635
rect 23447 67589 23525 67635
rect 23571 67589 23649 67635
rect 23695 67589 23773 67635
rect 23819 67589 23897 67635
rect 23943 67589 24021 67635
rect 24067 67589 24145 67635
rect 24191 67589 24269 67635
rect 24315 67589 24393 67635
rect 24439 67589 24517 67635
rect 24563 67589 24641 67635
rect 24687 67589 24765 67635
rect 24811 67589 24889 67635
rect 24935 67589 25013 67635
rect 25059 67589 25137 67635
rect 25183 67589 25261 67635
rect 25307 67589 25385 67635
rect 25431 67589 25509 67635
rect 25555 67589 25633 67635
rect 25679 67589 25757 67635
rect 25803 67589 25881 67635
rect 25927 67589 26005 67635
rect 26051 67589 26129 67635
rect 26175 67589 26253 67635
rect 26299 67589 26377 67635
rect 26423 67589 26501 67635
rect 26547 67589 26625 67635
rect 26671 67589 26749 67635
rect 26795 67589 26873 67635
rect 26919 67589 26997 67635
rect 27043 67589 27121 67635
rect 27167 67589 27245 67635
rect 27291 67589 27369 67635
rect 27415 67589 27493 67635
rect 27539 67589 27617 67635
rect 27663 67589 27741 67635
rect 27787 67589 27865 67635
rect 27911 67589 27989 67635
rect 28035 67589 28113 67635
rect 28159 67589 28237 67635
rect 28283 67589 28361 67635
rect 28407 67589 28485 67635
rect 28531 67589 28609 67635
rect 28655 67589 28733 67635
rect 28779 67589 28857 67635
rect 28903 67589 28981 67635
rect 29027 67589 29105 67635
rect 29151 67589 29229 67635
rect 29275 67589 29353 67635
rect 29399 67589 29477 67635
rect 29523 67589 29601 67635
rect 29647 67589 29725 67635
rect 29771 67589 29849 67635
rect 29895 67589 29973 67635
rect 30019 67589 30097 67635
rect 30143 67589 30221 67635
rect 30267 67589 30345 67635
rect 30391 67589 30469 67635
rect 30515 67589 30593 67635
rect 30639 67589 30717 67635
rect 30763 67589 30841 67635
rect 30887 67589 30965 67635
rect 31011 67589 31089 67635
rect 31135 67589 31213 67635
rect 31259 67589 31337 67635
rect 31383 67589 31461 67635
rect 31507 67589 31585 67635
rect 31631 67589 31709 67635
rect 31755 67589 31833 67635
rect 31879 67589 31957 67635
rect 32003 67589 32081 67635
rect 32127 67589 32205 67635
rect 32251 67589 32329 67635
rect 32375 67589 32453 67635
rect 32499 67589 32577 67635
rect 32623 67589 32701 67635
rect 32747 67589 32825 67635
rect 32871 67589 32949 67635
rect 32995 67589 33073 67635
rect 33119 67589 33197 67635
rect 33243 67589 33321 67635
rect 33367 67589 33445 67635
rect 33491 67589 33569 67635
rect 33615 67589 33693 67635
rect 33739 67589 33817 67635
rect 33863 67589 33941 67635
rect 33987 67589 34065 67635
rect 34111 67589 34189 67635
rect 34235 67589 34313 67635
rect 34359 67589 34437 67635
rect 34483 67589 34561 67635
rect 34607 67589 34685 67635
rect 34731 67589 34809 67635
rect 34855 67589 34933 67635
rect 34979 67589 35057 67635
rect 35103 67589 35181 67635
rect 35227 67589 35305 67635
rect 35351 67589 35429 67635
rect 35475 67589 35553 67635
rect 35599 67589 35677 67635
rect 35723 67589 35801 67635
rect 35847 67589 35925 67635
rect 35971 67589 36049 67635
rect 36095 67589 36173 67635
rect 36219 67589 36297 67635
rect 36343 67589 36421 67635
rect 36467 67589 36545 67635
rect 36591 67589 36669 67635
rect 36715 67589 36793 67635
rect 36839 67589 36917 67635
rect 36963 67589 37041 67635
rect 37087 67589 37165 67635
rect 37211 67589 37289 67635
rect 37335 67589 37413 67635
rect 37459 67589 37537 67635
rect 37583 67589 37661 67635
rect 37707 67589 37785 67635
rect 37831 67589 37909 67635
rect 37955 67589 38033 67635
rect 38079 67589 38157 67635
rect 38203 67589 38281 67635
rect 38327 67589 38405 67635
rect 38451 67589 38529 67635
rect 38575 67589 38653 67635
rect 38699 67589 38777 67635
rect 38823 67589 38901 67635
rect 38947 67589 39025 67635
rect 39071 67589 39149 67635
rect 39195 67589 39273 67635
rect 39319 67589 39397 67635
rect 39443 67589 39521 67635
rect 39567 67589 39645 67635
rect 39691 67589 39769 67635
rect 39815 67589 39893 67635
rect 39939 67589 40017 67635
rect 40063 67589 40141 67635
rect 40187 67589 40265 67635
rect 40311 67589 40389 67635
rect 40435 67589 40513 67635
rect 40559 67589 40637 67635
rect 40683 67589 40761 67635
rect 40807 67589 40885 67635
rect 40931 67589 41009 67635
rect 41055 67589 41133 67635
rect 41179 67589 41257 67635
rect 41303 67589 41381 67635
rect 41427 67589 41505 67635
rect 41551 67589 41629 67635
rect 41675 67589 41753 67635
rect 41799 67589 41877 67635
rect 41923 67589 42001 67635
rect 42047 67589 42125 67635
rect 42171 67589 42249 67635
rect 42295 67589 42373 67635
rect 42419 67589 42497 67635
rect 42543 67589 42621 67635
rect 42667 67589 42745 67635
rect 42791 67589 42869 67635
rect 42915 67589 42993 67635
rect 43039 67589 43117 67635
rect 43163 67589 43241 67635
rect 43287 67589 43365 67635
rect 43411 67589 43489 67635
rect 43535 67589 43613 67635
rect 43659 67589 43737 67635
rect 43783 67589 43861 67635
rect 43907 67589 43985 67635
rect 44031 67589 44109 67635
rect 44155 67589 44233 67635
rect 44279 67589 44357 67635
rect 44403 67589 44481 67635
rect 44527 67589 44605 67635
rect 44651 67589 44729 67635
rect 44775 67589 44853 67635
rect 44899 67589 44977 67635
rect 45023 67589 45101 67635
rect 45147 67589 45225 67635
rect 45271 67589 45349 67635
rect 45395 67589 45473 67635
rect 45519 67589 45597 67635
rect 45643 67589 45721 67635
rect 45767 67589 45845 67635
rect 45891 67589 45969 67635
rect 46015 67589 46093 67635
rect 46139 67589 46217 67635
rect 46263 67589 46341 67635
rect 46387 67589 46465 67635
rect 46511 67589 46589 67635
rect 46635 67589 46713 67635
rect 46759 67589 46837 67635
rect 46883 67589 46961 67635
rect 47007 67589 47085 67635
rect 47131 67589 47209 67635
rect 47255 67589 47333 67635
rect 47379 67589 47457 67635
rect 47503 67589 47581 67635
rect 47627 67589 47705 67635
rect 47751 67589 47829 67635
rect 47875 67589 47953 67635
rect 47999 67589 48077 67635
rect 48123 67589 48201 67635
rect 48247 67589 48325 67635
rect 48371 67589 48449 67635
rect 48495 67589 48573 67635
rect 48619 67589 48697 67635
rect 48743 67589 48821 67635
rect 48867 67589 48945 67635
rect 48991 67589 49069 67635
rect 49115 67589 49193 67635
rect 49239 67589 49317 67635
rect 49363 67589 49441 67635
rect 49487 67589 49565 67635
rect 49611 67589 49689 67635
rect 49735 67589 49813 67635
rect 49859 67589 49937 67635
rect 49983 67589 50061 67635
rect 50107 67589 50185 67635
rect 50231 67589 50309 67635
rect 50355 67589 50433 67635
rect 50479 67589 50557 67635
rect 50603 67589 50681 67635
rect 50727 67589 50805 67635
rect 50851 67589 50929 67635
rect 50975 67589 51053 67635
rect 51099 67589 51177 67635
rect 51223 67589 51301 67635
rect 51347 67589 51425 67635
rect 51471 67589 51549 67635
rect 51595 67589 51673 67635
rect 51719 67589 51797 67635
rect 51843 67589 51921 67635
rect 51967 67589 52045 67635
rect 52091 67589 52169 67635
rect 52215 67589 52293 67635
rect 52339 67589 52417 67635
rect 52463 67589 52541 67635
rect 52587 67589 52665 67635
rect 52711 67589 52789 67635
rect 52835 67589 52913 67635
rect 52959 67589 53037 67635
rect 53083 67589 53161 67635
rect 53207 67589 53285 67635
rect 53331 67589 53409 67635
rect 53455 67589 53533 67635
rect 53579 67589 53657 67635
rect 53703 67589 53781 67635
rect 53827 67589 53905 67635
rect 53951 67589 54029 67635
rect 54075 67589 54153 67635
rect 54199 67589 54277 67635
rect 54323 67589 54401 67635
rect 54447 67589 54525 67635
rect 54571 67589 54649 67635
rect 54695 67589 54773 67635
rect 54819 67589 54897 67635
rect 54943 67589 55021 67635
rect 55067 67589 55145 67635
rect 55191 67589 55269 67635
rect 55315 67589 55393 67635
rect 55439 67589 55517 67635
rect 55563 67589 55641 67635
rect 55687 67589 55765 67635
rect 55811 67589 55889 67635
rect 55935 67589 56013 67635
rect 56059 67589 56137 67635
rect 56183 67589 56261 67635
rect 56307 67589 56385 67635
rect 56431 67589 56509 67635
rect 56555 67589 56633 67635
rect 56679 67589 56757 67635
rect 56803 67589 56881 67635
rect 56927 67589 57005 67635
rect 57051 67589 57129 67635
rect 57175 67589 57253 67635
rect 57299 67589 57377 67635
rect 57423 67589 57501 67635
rect 57547 67589 57625 67635
rect 57671 67589 57749 67635
rect 57795 67589 57873 67635
rect 57919 67589 57997 67635
rect 58043 67589 58121 67635
rect 58167 67589 58245 67635
rect 58291 67589 58369 67635
rect 58415 67589 58493 67635
rect 58539 67589 58617 67635
rect 58663 67589 58741 67635
rect 58787 67589 58865 67635
rect 58911 67589 58989 67635
rect 59035 67589 59113 67635
rect 59159 67589 59237 67635
rect 59283 67589 59361 67635
rect 59407 67589 59485 67635
rect 59531 67589 59609 67635
rect 59655 67589 59733 67635
rect 59779 67589 59857 67635
rect 59903 67589 59981 67635
rect 60027 67589 60105 67635
rect 60151 67589 60229 67635
rect 60275 67589 60353 67635
rect 60399 67589 60477 67635
rect 60523 67589 60601 67635
rect 60647 67589 60725 67635
rect 60771 67589 60849 67635
rect 60895 67589 60973 67635
rect 61019 67589 61097 67635
rect 61143 67589 61221 67635
rect 61267 67589 61345 67635
rect 61391 67589 61469 67635
rect 61515 67589 61593 67635
rect 61639 67589 61717 67635
rect 61763 67589 61841 67635
rect 61887 67589 61965 67635
rect 62011 67589 62089 67635
rect 62135 67589 62213 67635
rect 62259 67589 62337 67635
rect 62383 67589 62461 67635
rect 62507 67589 62585 67635
rect 62631 67589 62709 67635
rect 62755 67589 62833 67635
rect 62879 67589 62957 67635
rect 63003 67589 63081 67635
rect 63127 67589 63205 67635
rect 63251 67589 63329 67635
rect 63375 67589 63453 67635
rect 63499 67589 63577 67635
rect 63623 67589 63701 67635
rect 63747 67589 63825 67635
rect 63871 67589 63949 67635
rect 63995 67589 64073 67635
rect 64119 67589 64197 67635
rect 64243 67589 64321 67635
rect 64367 67589 64445 67635
rect 64491 67589 64569 67635
rect 64615 67589 64693 67635
rect 64739 67589 64817 67635
rect 64863 67589 64941 67635
rect 64987 67589 65065 67635
rect 65111 67589 65189 67635
rect 65235 67589 65313 67635
rect 65359 67589 65437 67635
rect 65483 67589 65561 67635
rect 65607 67589 65685 67635
rect 65731 67589 65809 67635
rect 65855 67589 65933 67635
rect 65979 67589 66057 67635
rect 66103 67589 66181 67635
rect 66227 67589 66305 67635
rect 66351 67589 66429 67635
rect 66475 67589 66553 67635
rect 66599 67589 66677 67635
rect 66723 67589 66801 67635
rect 66847 67589 66925 67635
rect 66971 67589 67049 67635
rect 67095 67589 67173 67635
rect 67219 67589 67297 67635
rect 67343 67589 67421 67635
rect 67467 67589 67545 67635
rect 67591 67589 67669 67635
rect 67715 67589 67793 67635
rect 67839 67589 67917 67635
rect 67963 67589 68041 67635
rect 68087 67589 68165 67635
rect 68211 67589 68289 67635
rect 68335 67589 68413 67635
rect 68459 67589 68537 67635
rect 68583 67589 68661 67635
rect 68707 67589 68785 67635
rect 68831 67589 68909 67635
rect 68955 67589 69033 67635
rect 69079 67589 69157 67635
rect 69203 67589 69281 67635
rect 69327 67589 69405 67635
rect 69451 67589 69529 67635
rect 69575 67589 69653 67635
rect 69699 67589 69777 67635
rect 69823 67589 69901 67635
rect 69947 67589 70025 67635
rect 70071 67589 70149 67635
rect 70195 67589 70273 67635
rect 70319 67589 70397 67635
rect 70443 67589 70521 67635
rect 70567 67589 70645 67635
rect 70691 67589 70769 67635
rect 70815 67589 70893 67635
rect 70939 67589 71017 67635
rect 71063 67589 71141 67635
rect 71187 67589 71265 67635
rect 71311 67589 71389 67635
rect 71435 67589 71513 67635
rect 71559 67589 71637 67635
rect 71683 67589 71761 67635
rect 71807 67589 71885 67635
rect 71931 67589 72009 67635
rect 72055 67589 72133 67635
rect 72179 67589 72257 67635
rect 72303 67589 72381 67635
rect 72427 67589 72505 67635
rect 72551 67589 72629 67635
rect 72675 67589 72753 67635
rect 72799 67589 72877 67635
rect 72923 67589 73001 67635
rect 73047 67589 73125 67635
rect 73171 67589 73249 67635
rect 73295 67589 73373 67635
rect 73419 67589 73497 67635
rect 73543 67589 73621 67635
rect 73667 67589 73745 67635
rect 73791 67589 73869 67635
rect 73915 67589 73993 67635
rect 74039 67589 74117 67635
rect 74163 67589 74241 67635
rect 74287 67589 74365 67635
rect 74411 67589 74489 67635
rect 74535 67589 74613 67635
rect 74659 67589 74737 67635
rect 74783 67589 74861 67635
rect 74907 67589 74985 67635
rect 75031 67589 75109 67635
rect 75155 67589 75233 67635
rect 75279 67589 75357 67635
rect 75403 67589 75481 67635
rect 75527 67589 75605 67635
rect 75651 67589 75729 67635
rect 75775 67589 75853 67635
rect 75899 67589 75977 67635
rect 76023 67589 76101 67635
rect 76147 67589 76225 67635
rect 76271 67589 76349 67635
rect 76395 67589 76473 67635
rect 76519 67589 76597 67635
rect 76643 67589 76721 67635
rect 76767 67589 76845 67635
rect 76891 67589 76969 67635
rect 77015 67589 77093 67635
rect 77139 67589 77217 67635
rect 77263 67589 77341 67635
rect 77387 67589 77465 67635
rect 77511 67589 77589 67635
rect 77635 67589 77713 67635
rect 77759 67589 77837 67635
rect 77883 67589 77961 67635
rect 78007 67589 78085 67635
rect 78131 67589 78209 67635
rect 78255 67589 78333 67635
rect 78379 67589 78457 67635
rect 78503 67589 78581 67635
rect 78627 67589 78705 67635
rect 78751 67589 78829 67635
rect 78875 67589 78953 67635
rect 78999 67589 79077 67635
rect 79123 67589 79201 67635
rect 79247 67589 79325 67635
rect 79371 67589 79449 67635
rect 79495 67589 79573 67635
rect 79619 67589 79697 67635
rect 79743 67589 79821 67635
rect 79867 67589 79945 67635
rect 79991 67589 80069 67635
rect 80115 67589 80193 67635
rect 80239 67589 80317 67635
rect 80363 67589 80441 67635
rect 80487 67589 80565 67635
rect 80611 67589 80689 67635
rect 80735 67589 80813 67635
rect 80859 67589 80937 67635
rect 80983 67589 81061 67635
rect 81107 67589 81185 67635
rect 81231 67589 81309 67635
rect 81355 67589 81433 67635
rect 81479 67589 81557 67635
rect 81603 67589 81681 67635
rect 81727 67589 81805 67635
rect 81851 67589 81929 67635
rect 81975 67589 82053 67635
rect 82099 67589 82177 67635
rect 82223 67589 82301 67635
rect 82347 67589 82425 67635
rect 82471 67589 82549 67635
rect 82595 67589 82673 67635
rect 82719 67589 82797 67635
rect 82843 67589 82921 67635
rect 82967 67589 83045 67635
rect 83091 67589 83169 67635
rect 83215 67589 83293 67635
rect 83339 67589 83417 67635
rect 83463 67589 83541 67635
rect 83587 67589 83665 67635
rect 83711 67589 83789 67635
rect 83835 67589 83913 67635
rect 83959 67589 84037 67635
rect 84083 67589 84161 67635
rect 84207 67589 84285 67635
rect 84331 67589 84409 67635
rect 84455 67589 84533 67635
rect 84579 67589 84657 67635
rect 84703 67589 84781 67635
rect 84827 67589 84905 67635
rect 84951 67589 85029 67635
rect 85075 67589 85153 67635
rect 85199 67589 85277 67635
rect 85323 67589 85401 67635
rect 85447 67589 85525 67635
rect 85571 67589 85649 67635
rect 85695 67589 85816 67635
rect 70 67511 85816 67589
rect 70 67465 89 67511
rect 135 67465 213 67511
rect 259 67465 337 67511
rect 383 67465 461 67511
rect 507 67465 585 67511
rect 631 67465 709 67511
rect 755 67465 833 67511
rect 879 67465 957 67511
rect 1003 67465 1081 67511
rect 1127 67465 1205 67511
rect 1251 67465 1329 67511
rect 1375 67465 1453 67511
rect 1499 67465 1577 67511
rect 1623 67465 1701 67511
rect 1747 67465 1825 67511
rect 1871 67465 1949 67511
rect 1995 67465 2073 67511
rect 2119 67465 2197 67511
rect 2243 67465 2321 67511
rect 2367 67465 2445 67511
rect 2491 67465 2569 67511
rect 2615 67465 2693 67511
rect 2739 67465 2817 67511
rect 2863 67465 2941 67511
rect 2987 67465 3065 67511
rect 3111 67465 3189 67511
rect 3235 67465 3313 67511
rect 3359 67465 3437 67511
rect 3483 67465 3561 67511
rect 3607 67465 3685 67511
rect 3731 67465 3809 67511
rect 3855 67465 3933 67511
rect 3979 67465 4057 67511
rect 4103 67465 4181 67511
rect 4227 67465 4305 67511
rect 4351 67465 4429 67511
rect 4475 67465 4553 67511
rect 4599 67465 4677 67511
rect 4723 67465 4801 67511
rect 4847 67465 4925 67511
rect 4971 67465 5049 67511
rect 5095 67465 5173 67511
rect 5219 67465 5297 67511
rect 5343 67465 5421 67511
rect 5467 67465 5545 67511
rect 5591 67465 5669 67511
rect 5715 67465 5793 67511
rect 5839 67465 5917 67511
rect 5963 67465 6041 67511
rect 6087 67465 6165 67511
rect 6211 67465 6289 67511
rect 6335 67465 6413 67511
rect 6459 67465 6537 67511
rect 6583 67465 6661 67511
rect 6707 67465 6785 67511
rect 6831 67465 6909 67511
rect 6955 67465 7033 67511
rect 7079 67465 7157 67511
rect 7203 67465 7281 67511
rect 7327 67465 7405 67511
rect 7451 67465 7529 67511
rect 7575 67465 7653 67511
rect 7699 67465 7777 67511
rect 7823 67465 7901 67511
rect 7947 67465 8025 67511
rect 8071 67465 8149 67511
rect 8195 67465 8273 67511
rect 8319 67465 8397 67511
rect 8443 67465 8521 67511
rect 8567 67465 8645 67511
rect 8691 67465 8769 67511
rect 8815 67465 8893 67511
rect 8939 67465 9017 67511
rect 9063 67465 9141 67511
rect 9187 67465 9265 67511
rect 9311 67465 9389 67511
rect 9435 67465 9513 67511
rect 9559 67465 9637 67511
rect 9683 67465 9761 67511
rect 9807 67465 9885 67511
rect 9931 67465 10009 67511
rect 10055 67465 10133 67511
rect 10179 67465 10257 67511
rect 10303 67465 10381 67511
rect 10427 67465 10505 67511
rect 10551 67465 10629 67511
rect 10675 67465 10753 67511
rect 10799 67465 10877 67511
rect 10923 67465 11001 67511
rect 11047 67465 11125 67511
rect 11171 67465 11249 67511
rect 11295 67465 11373 67511
rect 11419 67465 11497 67511
rect 11543 67465 11621 67511
rect 11667 67465 11745 67511
rect 11791 67465 11869 67511
rect 11915 67465 11993 67511
rect 12039 67465 12117 67511
rect 12163 67465 12241 67511
rect 12287 67465 12365 67511
rect 12411 67465 12489 67511
rect 12535 67465 12613 67511
rect 12659 67465 12737 67511
rect 12783 67465 12861 67511
rect 12907 67465 12985 67511
rect 13031 67465 13109 67511
rect 13155 67465 13233 67511
rect 13279 67465 13357 67511
rect 13403 67465 13481 67511
rect 13527 67465 13605 67511
rect 13651 67465 13729 67511
rect 13775 67465 13853 67511
rect 13899 67465 13977 67511
rect 14023 67465 14101 67511
rect 14147 67465 14225 67511
rect 14271 67465 14349 67511
rect 14395 67465 14473 67511
rect 14519 67465 14597 67511
rect 14643 67465 14721 67511
rect 14767 67465 14845 67511
rect 14891 67465 14969 67511
rect 15015 67465 15093 67511
rect 15139 67465 15217 67511
rect 15263 67465 15341 67511
rect 15387 67465 15465 67511
rect 15511 67465 15589 67511
rect 15635 67465 15713 67511
rect 15759 67465 15837 67511
rect 15883 67465 15961 67511
rect 16007 67465 16085 67511
rect 16131 67465 16209 67511
rect 16255 67465 16333 67511
rect 16379 67465 16457 67511
rect 16503 67465 16581 67511
rect 16627 67465 16705 67511
rect 16751 67465 16829 67511
rect 16875 67465 16953 67511
rect 16999 67465 17077 67511
rect 17123 67465 17201 67511
rect 17247 67465 17325 67511
rect 17371 67465 17449 67511
rect 17495 67465 17573 67511
rect 17619 67465 17697 67511
rect 17743 67465 17821 67511
rect 17867 67465 17945 67511
rect 17991 67465 18069 67511
rect 18115 67465 18193 67511
rect 18239 67465 18317 67511
rect 18363 67465 18441 67511
rect 18487 67465 18565 67511
rect 18611 67465 18689 67511
rect 18735 67465 18813 67511
rect 18859 67465 18937 67511
rect 18983 67465 19061 67511
rect 19107 67465 19185 67511
rect 19231 67465 19309 67511
rect 19355 67465 19433 67511
rect 19479 67465 19557 67511
rect 19603 67465 19681 67511
rect 19727 67465 19805 67511
rect 19851 67465 19929 67511
rect 19975 67465 20053 67511
rect 20099 67465 20177 67511
rect 20223 67465 20301 67511
rect 20347 67465 20425 67511
rect 20471 67465 20549 67511
rect 20595 67465 20673 67511
rect 20719 67465 20797 67511
rect 20843 67465 20921 67511
rect 20967 67465 21045 67511
rect 21091 67465 21169 67511
rect 21215 67465 21293 67511
rect 21339 67465 21417 67511
rect 21463 67465 21541 67511
rect 21587 67465 21665 67511
rect 21711 67465 21789 67511
rect 21835 67465 21913 67511
rect 21959 67465 22037 67511
rect 22083 67465 22161 67511
rect 22207 67465 22285 67511
rect 22331 67465 22409 67511
rect 22455 67465 22533 67511
rect 22579 67465 22657 67511
rect 22703 67465 22781 67511
rect 22827 67465 22905 67511
rect 22951 67465 23029 67511
rect 23075 67465 23153 67511
rect 23199 67465 23277 67511
rect 23323 67465 23401 67511
rect 23447 67465 23525 67511
rect 23571 67465 23649 67511
rect 23695 67465 23773 67511
rect 23819 67465 23897 67511
rect 23943 67465 24021 67511
rect 24067 67465 24145 67511
rect 24191 67465 24269 67511
rect 24315 67465 24393 67511
rect 24439 67465 24517 67511
rect 24563 67465 24641 67511
rect 24687 67465 24765 67511
rect 24811 67465 24889 67511
rect 24935 67465 25013 67511
rect 25059 67465 25137 67511
rect 25183 67465 25261 67511
rect 25307 67465 25385 67511
rect 25431 67465 25509 67511
rect 25555 67465 25633 67511
rect 25679 67465 25757 67511
rect 25803 67465 25881 67511
rect 25927 67465 26005 67511
rect 26051 67465 26129 67511
rect 26175 67465 26253 67511
rect 26299 67465 26377 67511
rect 26423 67465 26501 67511
rect 26547 67465 26625 67511
rect 26671 67465 26749 67511
rect 26795 67465 26873 67511
rect 26919 67465 26997 67511
rect 27043 67465 27121 67511
rect 27167 67465 27245 67511
rect 27291 67465 27369 67511
rect 27415 67465 27493 67511
rect 27539 67465 27617 67511
rect 27663 67465 27741 67511
rect 27787 67465 27865 67511
rect 27911 67465 27989 67511
rect 28035 67465 28113 67511
rect 28159 67465 28237 67511
rect 28283 67465 28361 67511
rect 28407 67465 28485 67511
rect 28531 67465 28609 67511
rect 28655 67465 28733 67511
rect 28779 67465 28857 67511
rect 28903 67465 28981 67511
rect 29027 67465 29105 67511
rect 29151 67465 29229 67511
rect 29275 67465 29353 67511
rect 29399 67465 29477 67511
rect 29523 67465 29601 67511
rect 29647 67465 29725 67511
rect 29771 67465 29849 67511
rect 29895 67465 29973 67511
rect 30019 67465 30097 67511
rect 30143 67465 30221 67511
rect 30267 67465 30345 67511
rect 30391 67465 30469 67511
rect 30515 67465 30593 67511
rect 30639 67465 30717 67511
rect 30763 67465 30841 67511
rect 30887 67465 30965 67511
rect 31011 67465 31089 67511
rect 31135 67465 31213 67511
rect 31259 67465 31337 67511
rect 31383 67465 31461 67511
rect 31507 67465 31585 67511
rect 31631 67465 31709 67511
rect 31755 67465 31833 67511
rect 31879 67465 31957 67511
rect 32003 67465 32081 67511
rect 32127 67465 32205 67511
rect 32251 67465 32329 67511
rect 32375 67465 32453 67511
rect 32499 67465 32577 67511
rect 32623 67465 32701 67511
rect 32747 67465 32825 67511
rect 32871 67465 32949 67511
rect 32995 67465 33073 67511
rect 33119 67465 33197 67511
rect 33243 67465 33321 67511
rect 33367 67465 33445 67511
rect 33491 67465 33569 67511
rect 33615 67465 33693 67511
rect 33739 67465 33817 67511
rect 33863 67465 33941 67511
rect 33987 67465 34065 67511
rect 34111 67465 34189 67511
rect 34235 67465 34313 67511
rect 34359 67465 34437 67511
rect 34483 67465 34561 67511
rect 34607 67465 34685 67511
rect 34731 67465 34809 67511
rect 34855 67465 34933 67511
rect 34979 67465 35057 67511
rect 35103 67465 35181 67511
rect 35227 67465 35305 67511
rect 35351 67465 35429 67511
rect 35475 67465 35553 67511
rect 35599 67465 35677 67511
rect 35723 67465 35801 67511
rect 35847 67465 35925 67511
rect 35971 67465 36049 67511
rect 36095 67465 36173 67511
rect 36219 67465 36297 67511
rect 36343 67465 36421 67511
rect 36467 67465 36545 67511
rect 36591 67465 36669 67511
rect 36715 67465 36793 67511
rect 36839 67465 36917 67511
rect 36963 67465 37041 67511
rect 37087 67465 37165 67511
rect 37211 67465 37289 67511
rect 37335 67465 37413 67511
rect 37459 67465 37537 67511
rect 37583 67465 37661 67511
rect 37707 67465 37785 67511
rect 37831 67465 37909 67511
rect 37955 67465 38033 67511
rect 38079 67465 38157 67511
rect 38203 67465 38281 67511
rect 38327 67465 38405 67511
rect 38451 67465 38529 67511
rect 38575 67465 38653 67511
rect 38699 67465 38777 67511
rect 38823 67465 38901 67511
rect 38947 67465 39025 67511
rect 39071 67465 39149 67511
rect 39195 67465 39273 67511
rect 39319 67465 39397 67511
rect 39443 67465 39521 67511
rect 39567 67465 39645 67511
rect 39691 67465 39769 67511
rect 39815 67465 39893 67511
rect 39939 67465 40017 67511
rect 40063 67465 40141 67511
rect 40187 67465 40265 67511
rect 40311 67465 40389 67511
rect 40435 67465 40513 67511
rect 40559 67465 40637 67511
rect 40683 67465 40761 67511
rect 40807 67465 40885 67511
rect 40931 67465 41009 67511
rect 41055 67465 41133 67511
rect 41179 67465 41257 67511
rect 41303 67465 41381 67511
rect 41427 67465 41505 67511
rect 41551 67465 41629 67511
rect 41675 67465 41753 67511
rect 41799 67465 41877 67511
rect 41923 67465 42001 67511
rect 42047 67465 42125 67511
rect 42171 67465 42249 67511
rect 42295 67465 42373 67511
rect 42419 67465 42497 67511
rect 42543 67465 42621 67511
rect 42667 67465 42745 67511
rect 42791 67465 42869 67511
rect 42915 67465 42993 67511
rect 43039 67465 43117 67511
rect 43163 67465 43241 67511
rect 43287 67465 43365 67511
rect 43411 67465 43489 67511
rect 43535 67465 43613 67511
rect 43659 67465 43737 67511
rect 43783 67465 43861 67511
rect 43907 67465 43985 67511
rect 44031 67465 44109 67511
rect 44155 67465 44233 67511
rect 44279 67465 44357 67511
rect 44403 67465 44481 67511
rect 44527 67465 44605 67511
rect 44651 67465 44729 67511
rect 44775 67465 44853 67511
rect 44899 67465 44977 67511
rect 45023 67465 45101 67511
rect 45147 67465 45225 67511
rect 45271 67465 45349 67511
rect 45395 67465 45473 67511
rect 45519 67465 45597 67511
rect 45643 67465 45721 67511
rect 45767 67465 45845 67511
rect 45891 67465 45969 67511
rect 46015 67465 46093 67511
rect 46139 67465 46217 67511
rect 46263 67465 46341 67511
rect 46387 67465 46465 67511
rect 46511 67465 46589 67511
rect 46635 67465 46713 67511
rect 46759 67465 46837 67511
rect 46883 67465 46961 67511
rect 47007 67465 47085 67511
rect 47131 67465 47209 67511
rect 47255 67465 47333 67511
rect 47379 67465 47457 67511
rect 47503 67465 47581 67511
rect 47627 67465 47705 67511
rect 47751 67465 47829 67511
rect 47875 67465 47953 67511
rect 47999 67465 48077 67511
rect 48123 67465 48201 67511
rect 48247 67465 48325 67511
rect 48371 67465 48449 67511
rect 48495 67465 48573 67511
rect 48619 67465 48697 67511
rect 48743 67465 48821 67511
rect 48867 67465 48945 67511
rect 48991 67465 49069 67511
rect 49115 67465 49193 67511
rect 49239 67465 49317 67511
rect 49363 67465 49441 67511
rect 49487 67465 49565 67511
rect 49611 67465 49689 67511
rect 49735 67465 49813 67511
rect 49859 67465 49937 67511
rect 49983 67465 50061 67511
rect 50107 67465 50185 67511
rect 50231 67465 50309 67511
rect 50355 67465 50433 67511
rect 50479 67465 50557 67511
rect 50603 67465 50681 67511
rect 50727 67465 50805 67511
rect 50851 67465 50929 67511
rect 50975 67465 51053 67511
rect 51099 67465 51177 67511
rect 51223 67465 51301 67511
rect 51347 67465 51425 67511
rect 51471 67465 51549 67511
rect 51595 67465 51673 67511
rect 51719 67465 51797 67511
rect 51843 67465 51921 67511
rect 51967 67465 52045 67511
rect 52091 67465 52169 67511
rect 52215 67465 52293 67511
rect 52339 67465 52417 67511
rect 52463 67465 52541 67511
rect 52587 67465 52665 67511
rect 52711 67465 52789 67511
rect 52835 67465 52913 67511
rect 52959 67465 53037 67511
rect 53083 67465 53161 67511
rect 53207 67465 53285 67511
rect 53331 67465 53409 67511
rect 53455 67465 53533 67511
rect 53579 67465 53657 67511
rect 53703 67465 53781 67511
rect 53827 67465 53905 67511
rect 53951 67465 54029 67511
rect 54075 67465 54153 67511
rect 54199 67465 54277 67511
rect 54323 67465 54401 67511
rect 54447 67465 54525 67511
rect 54571 67465 54649 67511
rect 54695 67465 54773 67511
rect 54819 67465 54897 67511
rect 54943 67465 55021 67511
rect 55067 67465 55145 67511
rect 55191 67465 55269 67511
rect 55315 67465 55393 67511
rect 55439 67465 55517 67511
rect 55563 67465 55641 67511
rect 55687 67465 55765 67511
rect 55811 67465 55889 67511
rect 55935 67465 56013 67511
rect 56059 67465 56137 67511
rect 56183 67465 56261 67511
rect 56307 67465 56385 67511
rect 56431 67465 56509 67511
rect 56555 67465 56633 67511
rect 56679 67465 56757 67511
rect 56803 67465 56881 67511
rect 56927 67465 57005 67511
rect 57051 67465 57129 67511
rect 57175 67465 57253 67511
rect 57299 67465 57377 67511
rect 57423 67465 57501 67511
rect 57547 67465 57625 67511
rect 57671 67465 57749 67511
rect 57795 67465 57873 67511
rect 57919 67465 57997 67511
rect 58043 67465 58121 67511
rect 58167 67465 58245 67511
rect 58291 67465 58369 67511
rect 58415 67465 58493 67511
rect 58539 67465 58617 67511
rect 58663 67465 58741 67511
rect 58787 67465 58865 67511
rect 58911 67465 58989 67511
rect 59035 67465 59113 67511
rect 59159 67465 59237 67511
rect 59283 67465 59361 67511
rect 59407 67465 59485 67511
rect 59531 67465 59609 67511
rect 59655 67465 59733 67511
rect 59779 67465 59857 67511
rect 59903 67465 59981 67511
rect 60027 67465 60105 67511
rect 60151 67465 60229 67511
rect 60275 67465 60353 67511
rect 60399 67465 60477 67511
rect 60523 67465 60601 67511
rect 60647 67465 60725 67511
rect 60771 67465 60849 67511
rect 60895 67465 60973 67511
rect 61019 67465 61097 67511
rect 61143 67465 61221 67511
rect 61267 67465 61345 67511
rect 61391 67465 61469 67511
rect 61515 67465 61593 67511
rect 61639 67465 61717 67511
rect 61763 67465 61841 67511
rect 61887 67465 61965 67511
rect 62011 67465 62089 67511
rect 62135 67465 62213 67511
rect 62259 67465 62337 67511
rect 62383 67465 62461 67511
rect 62507 67465 62585 67511
rect 62631 67465 62709 67511
rect 62755 67465 62833 67511
rect 62879 67465 62957 67511
rect 63003 67465 63081 67511
rect 63127 67465 63205 67511
rect 63251 67465 63329 67511
rect 63375 67465 63453 67511
rect 63499 67465 63577 67511
rect 63623 67465 63701 67511
rect 63747 67465 63825 67511
rect 63871 67465 63949 67511
rect 63995 67465 64073 67511
rect 64119 67465 64197 67511
rect 64243 67465 64321 67511
rect 64367 67465 64445 67511
rect 64491 67465 64569 67511
rect 64615 67465 64693 67511
rect 64739 67465 64817 67511
rect 64863 67465 64941 67511
rect 64987 67465 65065 67511
rect 65111 67465 65189 67511
rect 65235 67465 65313 67511
rect 65359 67465 65437 67511
rect 65483 67465 65561 67511
rect 65607 67465 65685 67511
rect 65731 67465 65809 67511
rect 65855 67465 65933 67511
rect 65979 67465 66057 67511
rect 66103 67465 66181 67511
rect 66227 67465 66305 67511
rect 66351 67465 66429 67511
rect 66475 67465 66553 67511
rect 66599 67465 66677 67511
rect 66723 67465 66801 67511
rect 66847 67465 66925 67511
rect 66971 67465 67049 67511
rect 67095 67465 67173 67511
rect 67219 67465 67297 67511
rect 67343 67465 67421 67511
rect 67467 67465 67545 67511
rect 67591 67465 67669 67511
rect 67715 67465 67793 67511
rect 67839 67465 67917 67511
rect 67963 67465 68041 67511
rect 68087 67465 68165 67511
rect 68211 67465 68289 67511
rect 68335 67465 68413 67511
rect 68459 67465 68537 67511
rect 68583 67465 68661 67511
rect 68707 67465 68785 67511
rect 68831 67465 68909 67511
rect 68955 67465 69033 67511
rect 69079 67465 69157 67511
rect 69203 67465 69281 67511
rect 69327 67465 69405 67511
rect 69451 67465 69529 67511
rect 69575 67465 69653 67511
rect 69699 67465 69777 67511
rect 69823 67465 69901 67511
rect 69947 67465 70025 67511
rect 70071 67465 70149 67511
rect 70195 67465 70273 67511
rect 70319 67465 70397 67511
rect 70443 67465 70521 67511
rect 70567 67465 70645 67511
rect 70691 67465 70769 67511
rect 70815 67465 70893 67511
rect 70939 67465 71017 67511
rect 71063 67465 71141 67511
rect 71187 67465 71265 67511
rect 71311 67465 71389 67511
rect 71435 67465 71513 67511
rect 71559 67465 71637 67511
rect 71683 67465 71761 67511
rect 71807 67465 71885 67511
rect 71931 67465 72009 67511
rect 72055 67465 72133 67511
rect 72179 67465 72257 67511
rect 72303 67465 72381 67511
rect 72427 67465 72505 67511
rect 72551 67465 72629 67511
rect 72675 67465 72753 67511
rect 72799 67465 72877 67511
rect 72923 67465 73001 67511
rect 73047 67465 73125 67511
rect 73171 67465 73249 67511
rect 73295 67465 73373 67511
rect 73419 67465 73497 67511
rect 73543 67465 73621 67511
rect 73667 67465 73745 67511
rect 73791 67465 73869 67511
rect 73915 67465 73993 67511
rect 74039 67465 74117 67511
rect 74163 67465 74241 67511
rect 74287 67465 74365 67511
rect 74411 67465 74489 67511
rect 74535 67465 74613 67511
rect 74659 67465 74737 67511
rect 74783 67465 74861 67511
rect 74907 67465 74985 67511
rect 75031 67465 75109 67511
rect 75155 67465 75233 67511
rect 75279 67465 75357 67511
rect 75403 67465 75481 67511
rect 75527 67465 75605 67511
rect 75651 67465 75729 67511
rect 75775 67465 75853 67511
rect 75899 67465 75977 67511
rect 76023 67465 76101 67511
rect 76147 67465 76225 67511
rect 76271 67465 76349 67511
rect 76395 67465 76473 67511
rect 76519 67465 76597 67511
rect 76643 67465 76721 67511
rect 76767 67465 76845 67511
rect 76891 67465 76969 67511
rect 77015 67465 77093 67511
rect 77139 67465 77217 67511
rect 77263 67465 77341 67511
rect 77387 67465 77465 67511
rect 77511 67465 77589 67511
rect 77635 67465 77713 67511
rect 77759 67465 77837 67511
rect 77883 67465 77961 67511
rect 78007 67465 78085 67511
rect 78131 67465 78209 67511
rect 78255 67465 78333 67511
rect 78379 67465 78457 67511
rect 78503 67465 78581 67511
rect 78627 67465 78705 67511
rect 78751 67465 78829 67511
rect 78875 67465 78953 67511
rect 78999 67465 79077 67511
rect 79123 67465 79201 67511
rect 79247 67465 79325 67511
rect 79371 67465 79449 67511
rect 79495 67465 79573 67511
rect 79619 67465 79697 67511
rect 79743 67465 79821 67511
rect 79867 67465 79945 67511
rect 79991 67465 80069 67511
rect 80115 67465 80193 67511
rect 80239 67465 80317 67511
rect 80363 67465 80441 67511
rect 80487 67465 80565 67511
rect 80611 67465 80689 67511
rect 80735 67465 80813 67511
rect 80859 67465 80937 67511
rect 80983 67465 81061 67511
rect 81107 67465 81185 67511
rect 81231 67465 81309 67511
rect 81355 67465 81433 67511
rect 81479 67465 81557 67511
rect 81603 67465 81681 67511
rect 81727 67465 81805 67511
rect 81851 67465 81929 67511
rect 81975 67465 82053 67511
rect 82099 67465 82177 67511
rect 82223 67465 82301 67511
rect 82347 67465 82425 67511
rect 82471 67465 82549 67511
rect 82595 67465 82673 67511
rect 82719 67465 82797 67511
rect 82843 67465 82921 67511
rect 82967 67465 83045 67511
rect 83091 67465 83169 67511
rect 83215 67465 83293 67511
rect 83339 67465 83417 67511
rect 83463 67465 83541 67511
rect 83587 67465 83665 67511
rect 83711 67465 83789 67511
rect 83835 67465 83913 67511
rect 83959 67465 84037 67511
rect 84083 67465 84161 67511
rect 84207 67465 84285 67511
rect 84331 67465 84409 67511
rect 84455 67465 84533 67511
rect 84579 67465 84657 67511
rect 84703 67465 84781 67511
rect 84827 67465 84905 67511
rect 84951 67465 85029 67511
rect 85075 67465 85153 67511
rect 85199 67465 85277 67511
rect 85323 67465 85401 67511
rect 85447 67465 85525 67511
rect 85571 67465 85649 67511
rect 85695 67465 85816 67511
rect 70 67446 85816 67465
rect 70 67363 454 67446
rect 70 1117 89 67363
rect 435 1117 454 67363
rect 70 1034 454 1117
rect 27097 67363 27481 67382
rect 27097 1117 27116 67363
rect 27462 1117 27481 67363
rect 57005 67363 57389 67382
rect 27545 67342 28429 67361
rect 27545 35996 27564 67342
rect 28410 35996 28429 67342
rect 27545 35977 28429 35996
rect 56091 67342 56975 67361
rect 56091 35996 56110 67342
rect 56956 35996 56975 67342
rect 56091 35977 56975 35996
rect 27545 34588 56929 34607
rect 27545 34242 27564 34588
rect 56910 34242 56929 34588
rect 27545 34223 56929 34242
rect 27097 1034 27481 1117
rect 57005 1117 57024 67363
rect 57370 1117 57389 67363
rect 57005 1034 57389 1117
rect 85432 67363 85816 67446
rect 85432 1117 85451 67363
rect 85797 1117 85816 67363
rect 85432 1034 85816 1117
rect 70 1015 85816 1034
rect 70 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85816 1015
rect 70 891 85816 969
rect 70 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85816 891
rect 70 767 85816 845
rect 70 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85816 767
rect 70 643 85816 721
rect 70 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85816 643
rect 70 578 85816 597
<< psubdiffcont >>
rect 89 67837 135 67883
rect 213 67837 259 67883
rect 337 67837 383 67883
rect 461 67837 507 67883
rect 585 67837 631 67883
rect 709 67837 755 67883
rect 833 67837 879 67883
rect 957 67837 1003 67883
rect 1081 67837 1127 67883
rect 1205 67837 1251 67883
rect 1329 67837 1375 67883
rect 1453 67837 1499 67883
rect 1577 67837 1623 67883
rect 1701 67837 1747 67883
rect 1825 67837 1871 67883
rect 1949 67837 1995 67883
rect 2073 67837 2119 67883
rect 2197 67837 2243 67883
rect 2321 67837 2367 67883
rect 2445 67837 2491 67883
rect 2569 67837 2615 67883
rect 2693 67837 2739 67883
rect 2817 67837 2863 67883
rect 2941 67837 2987 67883
rect 3065 67837 3111 67883
rect 3189 67837 3235 67883
rect 3313 67837 3359 67883
rect 3437 67837 3483 67883
rect 3561 67837 3607 67883
rect 3685 67837 3731 67883
rect 3809 67837 3855 67883
rect 3933 67837 3979 67883
rect 4057 67837 4103 67883
rect 4181 67837 4227 67883
rect 4305 67837 4351 67883
rect 4429 67837 4475 67883
rect 4553 67837 4599 67883
rect 4677 67837 4723 67883
rect 4801 67837 4847 67883
rect 4925 67837 4971 67883
rect 5049 67837 5095 67883
rect 5173 67837 5219 67883
rect 5297 67837 5343 67883
rect 5421 67837 5467 67883
rect 5545 67837 5591 67883
rect 5669 67837 5715 67883
rect 5793 67837 5839 67883
rect 5917 67837 5963 67883
rect 6041 67837 6087 67883
rect 6165 67837 6211 67883
rect 6289 67837 6335 67883
rect 6413 67837 6459 67883
rect 6537 67837 6583 67883
rect 6661 67837 6707 67883
rect 6785 67837 6831 67883
rect 6909 67837 6955 67883
rect 7033 67837 7079 67883
rect 7157 67837 7203 67883
rect 7281 67837 7327 67883
rect 7405 67837 7451 67883
rect 7529 67837 7575 67883
rect 7653 67837 7699 67883
rect 7777 67837 7823 67883
rect 7901 67837 7947 67883
rect 8025 67837 8071 67883
rect 8149 67837 8195 67883
rect 8273 67837 8319 67883
rect 8397 67837 8443 67883
rect 8521 67837 8567 67883
rect 8645 67837 8691 67883
rect 8769 67837 8815 67883
rect 8893 67837 8939 67883
rect 9017 67837 9063 67883
rect 9141 67837 9187 67883
rect 9265 67837 9311 67883
rect 9389 67837 9435 67883
rect 9513 67837 9559 67883
rect 9637 67837 9683 67883
rect 9761 67837 9807 67883
rect 9885 67837 9931 67883
rect 10009 67837 10055 67883
rect 10133 67837 10179 67883
rect 10257 67837 10303 67883
rect 10381 67837 10427 67883
rect 10505 67837 10551 67883
rect 10629 67837 10675 67883
rect 10753 67837 10799 67883
rect 10877 67837 10923 67883
rect 11001 67837 11047 67883
rect 11125 67837 11171 67883
rect 11249 67837 11295 67883
rect 11373 67837 11419 67883
rect 11497 67837 11543 67883
rect 11621 67837 11667 67883
rect 11745 67837 11791 67883
rect 11869 67837 11915 67883
rect 11993 67837 12039 67883
rect 12117 67837 12163 67883
rect 12241 67837 12287 67883
rect 12365 67837 12411 67883
rect 12489 67837 12535 67883
rect 12613 67837 12659 67883
rect 12737 67837 12783 67883
rect 12861 67837 12907 67883
rect 12985 67837 13031 67883
rect 13109 67837 13155 67883
rect 13233 67837 13279 67883
rect 13357 67837 13403 67883
rect 13481 67837 13527 67883
rect 13605 67837 13651 67883
rect 13729 67837 13775 67883
rect 13853 67837 13899 67883
rect 13977 67837 14023 67883
rect 14101 67837 14147 67883
rect 14225 67837 14271 67883
rect 14349 67837 14395 67883
rect 14473 67837 14519 67883
rect 14597 67837 14643 67883
rect 14721 67837 14767 67883
rect 14845 67837 14891 67883
rect 14969 67837 15015 67883
rect 15093 67837 15139 67883
rect 15217 67837 15263 67883
rect 15341 67837 15387 67883
rect 15465 67837 15511 67883
rect 15589 67837 15635 67883
rect 15713 67837 15759 67883
rect 15837 67837 15883 67883
rect 15961 67837 16007 67883
rect 16085 67837 16131 67883
rect 16209 67837 16255 67883
rect 16333 67837 16379 67883
rect 16457 67837 16503 67883
rect 16581 67837 16627 67883
rect 16705 67837 16751 67883
rect 16829 67837 16875 67883
rect 16953 67837 16999 67883
rect 17077 67837 17123 67883
rect 17201 67837 17247 67883
rect 17325 67837 17371 67883
rect 17449 67837 17495 67883
rect 17573 67837 17619 67883
rect 17697 67837 17743 67883
rect 17821 67837 17867 67883
rect 17945 67837 17991 67883
rect 18069 67837 18115 67883
rect 18193 67837 18239 67883
rect 18317 67837 18363 67883
rect 18441 67837 18487 67883
rect 18565 67837 18611 67883
rect 18689 67837 18735 67883
rect 18813 67837 18859 67883
rect 18937 67837 18983 67883
rect 19061 67837 19107 67883
rect 19185 67837 19231 67883
rect 19309 67837 19355 67883
rect 19433 67837 19479 67883
rect 19557 67837 19603 67883
rect 19681 67837 19727 67883
rect 19805 67837 19851 67883
rect 19929 67837 19975 67883
rect 20053 67837 20099 67883
rect 20177 67837 20223 67883
rect 20301 67837 20347 67883
rect 20425 67837 20471 67883
rect 20549 67837 20595 67883
rect 20673 67837 20719 67883
rect 20797 67837 20843 67883
rect 20921 67837 20967 67883
rect 21045 67837 21091 67883
rect 21169 67837 21215 67883
rect 21293 67837 21339 67883
rect 21417 67837 21463 67883
rect 21541 67837 21587 67883
rect 21665 67837 21711 67883
rect 21789 67837 21835 67883
rect 21913 67837 21959 67883
rect 22037 67837 22083 67883
rect 22161 67837 22207 67883
rect 22285 67837 22331 67883
rect 22409 67837 22455 67883
rect 22533 67837 22579 67883
rect 22657 67837 22703 67883
rect 22781 67837 22827 67883
rect 22905 67837 22951 67883
rect 23029 67837 23075 67883
rect 23153 67837 23199 67883
rect 23277 67837 23323 67883
rect 23401 67837 23447 67883
rect 23525 67837 23571 67883
rect 23649 67837 23695 67883
rect 23773 67837 23819 67883
rect 23897 67837 23943 67883
rect 24021 67837 24067 67883
rect 24145 67837 24191 67883
rect 24269 67837 24315 67883
rect 24393 67837 24439 67883
rect 24517 67837 24563 67883
rect 24641 67837 24687 67883
rect 24765 67837 24811 67883
rect 24889 67837 24935 67883
rect 25013 67837 25059 67883
rect 25137 67837 25183 67883
rect 25261 67837 25307 67883
rect 25385 67837 25431 67883
rect 25509 67837 25555 67883
rect 25633 67837 25679 67883
rect 25757 67837 25803 67883
rect 25881 67837 25927 67883
rect 26005 67837 26051 67883
rect 26129 67837 26175 67883
rect 26253 67837 26299 67883
rect 26377 67837 26423 67883
rect 26501 67837 26547 67883
rect 26625 67837 26671 67883
rect 26749 67837 26795 67883
rect 26873 67837 26919 67883
rect 26997 67837 27043 67883
rect 27121 67837 27167 67883
rect 27245 67837 27291 67883
rect 27369 67837 27415 67883
rect 27493 67837 27539 67883
rect 27617 67837 27663 67883
rect 27741 67837 27787 67883
rect 27865 67837 27911 67883
rect 27989 67837 28035 67883
rect 28113 67837 28159 67883
rect 28237 67837 28283 67883
rect 28361 67837 28407 67883
rect 28485 67837 28531 67883
rect 28609 67837 28655 67883
rect 28733 67837 28779 67883
rect 28857 67837 28903 67883
rect 28981 67837 29027 67883
rect 29105 67837 29151 67883
rect 29229 67837 29275 67883
rect 29353 67837 29399 67883
rect 29477 67837 29523 67883
rect 29601 67837 29647 67883
rect 29725 67837 29771 67883
rect 29849 67837 29895 67883
rect 29973 67837 30019 67883
rect 30097 67837 30143 67883
rect 30221 67837 30267 67883
rect 30345 67837 30391 67883
rect 30469 67837 30515 67883
rect 30593 67837 30639 67883
rect 30717 67837 30763 67883
rect 30841 67837 30887 67883
rect 30965 67837 31011 67883
rect 31089 67837 31135 67883
rect 31213 67837 31259 67883
rect 31337 67837 31383 67883
rect 31461 67837 31507 67883
rect 31585 67837 31631 67883
rect 31709 67837 31755 67883
rect 31833 67837 31879 67883
rect 31957 67837 32003 67883
rect 32081 67837 32127 67883
rect 32205 67837 32251 67883
rect 32329 67837 32375 67883
rect 32453 67837 32499 67883
rect 32577 67837 32623 67883
rect 32701 67837 32747 67883
rect 32825 67837 32871 67883
rect 32949 67837 32995 67883
rect 33073 67837 33119 67883
rect 33197 67837 33243 67883
rect 33321 67837 33367 67883
rect 33445 67837 33491 67883
rect 33569 67837 33615 67883
rect 33693 67837 33739 67883
rect 33817 67837 33863 67883
rect 33941 67837 33987 67883
rect 34065 67837 34111 67883
rect 34189 67837 34235 67883
rect 34313 67837 34359 67883
rect 34437 67837 34483 67883
rect 34561 67837 34607 67883
rect 34685 67837 34731 67883
rect 34809 67837 34855 67883
rect 34933 67837 34979 67883
rect 35057 67837 35103 67883
rect 35181 67837 35227 67883
rect 35305 67837 35351 67883
rect 35429 67837 35475 67883
rect 35553 67837 35599 67883
rect 35677 67837 35723 67883
rect 35801 67837 35847 67883
rect 35925 67837 35971 67883
rect 36049 67837 36095 67883
rect 36173 67837 36219 67883
rect 36297 67837 36343 67883
rect 36421 67837 36467 67883
rect 36545 67837 36591 67883
rect 36669 67837 36715 67883
rect 36793 67837 36839 67883
rect 36917 67837 36963 67883
rect 37041 67837 37087 67883
rect 37165 67837 37211 67883
rect 37289 67837 37335 67883
rect 37413 67837 37459 67883
rect 37537 67837 37583 67883
rect 37661 67837 37707 67883
rect 37785 67837 37831 67883
rect 37909 67837 37955 67883
rect 38033 67837 38079 67883
rect 38157 67837 38203 67883
rect 38281 67837 38327 67883
rect 38405 67837 38451 67883
rect 38529 67837 38575 67883
rect 38653 67837 38699 67883
rect 38777 67837 38823 67883
rect 38901 67837 38947 67883
rect 39025 67837 39071 67883
rect 39149 67837 39195 67883
rect 39273 67837 39319 67883
rect 39397 67837 39443 67883
rect 39521 67837 39567 67883
rect 39645 67837 39691 67883
rect 39769 67837 39815 67883
rect 39893 67837 39939 67883
rect 40017 67837 40063 67883
rect 40141 67837 40187 67883
rect 40265 67837 40311 67883
rect 40389 67837 40435 67883
rect 40513 67837 40559 67883
rect 40637 67837 40683 67883
rect 40761 67837 40807 67883
rect 40885 67837 40931 67883
rect 41009 67837 41055 67883
rect 41133 67837 41179 67883
rect 41257 67837 41303 67883
rect 41381 67837 41427 67883
rect 41505 67837 41551 67883
rect 41629 67837 41675 67883
rect 41753 67837 41799 67883
rect 41877 67837 41923 67883
rect 42001 67837 42047 67883
rect 42125 67837 42171 67883
rect 42249 67837 42295 67883
rect 42373 67837 42419 67883
rect 42497 67837 42543 67883
rect 42621 67837 42667 67883
rect 42745 67837 42791 67883
rect 42869 67837 42915 67883
rect 42993 67837 43039 67883
rect 43117 67837 43163 67883
rect 43241 67837 43287 67883
rect 43365 67837 43411 67883
rect 43489 67837 43535 67883
rect 43613 67837 43659 67883
rect 43737 67837 43783 67883
rect 43861 67837 43907 67883
rect 43985 67837 44031 67883
rect 44109 67837 44155 67883
rect 44233 67837 44279 67883
rect 44357 67837 44403 67883
rect 44481 67837 44527 67883
rect 44605 67837 44651 67883
rect 44729 67837 44775 67883
rect 44853 67837 44899 67883
rect 44977 67837 45023 67883
rect 45101 67837 45147 67883
rect 45225 67837 45271 67883
rect 45349 67837 45395 67883
rect 45473 67837 45519 67883
rect 45597 67837 45643 67883
rect 45721 67837 45767 67883
rect 45845 67837 45891 67883
rect 45969 67837 46015 67883
rect 46093 67837 46139 67883
rect 46217 67837 46263 67883
rect 46341 67837 46387 67883
rect 46465 67837 46511 67883
rect 46589 67837 46635 67883
rect 46713 67837 46759 67883
rect 46837 67837 46883 67883
rect 46961 67837 47007 67883
rect 47085 67837 47131 67883
rect 47209 67837 47255 67883
rect 47333 67837 47379 67883
rect 47457 67837 47503 67883
rect 47581 67837 47627 67883
rect 47705 67837 47751 67883
rect 47829 67837 47875 67883
rect 47953 67837 47999 67883
rect 48077 67837 48123 67883
rect 48201 67837 48247 67883
rect 48325 67837 48371 67883
rect 48449 67837 48495 67883
rect 48573 67837 48619 67883
rect 48697 67837 48743 67883
rect 48821 67837 48867 67883
rect 48945 67837 48991 67883
rect 49069 67837 49115 67883
rect 49193 67837 49239 67883
rect 49317 67837 49363 67883
rect 49441 67837 49487 67883
rect 49565 67837 49611 67883
rect 49689 67837 49735 67883
rect 49813 67837 49859 67883
rect 49937 67837 49983 67883
rect 50061 67837 50107 67883
rect 50185 67837 50231 67883
rect 50309 67837 50355 67883
rect 50433 67837 50479 67883
rect 50557 67837 50603 67883
rect 50681 67837 50727 67883
rect 50805 67837 50851 67883
rect 50929 67837 50975 67883
rect 51053 67837 51099 67883
rect 51177 67837 51223 67883
rect 51301 67837 51347 67883
rect 51425 67837 51471 67883
rect 51549 67837 51595 67883
rect 51673 67837 51719 67883
rect 51797 67837 51843 67883
rect 51921 67837 51967 67883
rect 52045 67837 52091 67883
rect 52169 67837 52215 67883
rect 52293 67837 52339 67883
rect 52417 67837 52463 67883
rect 52541 67837 52587 67883
rect 52665 67837 52711 67883
rect 52789 67837 52835 67883
rect 52913 67837 52959 67883
rect 53037 67837 53083 67883
rect 53161 67837 53207 67883
rect 53285 67837 53331 67883
rect 53409 67837 53455 67883
rect 53533 67837 53579 67883
rect 53657 67837 53703 67883
rect 53781 67837 53827 67883
rect 53905 67837 53951 67883
rect 54029 67837 54075 67883
rect 54153 67837 54199 67883
rect 54277 67837 54323 67883
rect 54401 67837 54447 67883
rect 54525 67837 54571 67883
rect 54649 67837 54695 67883
rect 54773 67837 54819 67883
rect 54897 67837 54943 67883
rect 55021 67837 55067 67883
rect 55145 67837 55191 67883
rect 55269 67837 55315 67883
rect 55393 67837 55439 67883
rect 55517 67837 55563 67883
rect 55641 67837 55687 67883
rect 55765 67837 55811 67883
rect 55889 67837 55935 67883
rect 56013 67837 56059 67883
rect 56137 67837 56183 67883
rect 56261 67837 56307 67883
rect 56385 67837 56431 67883
rect 56509 67837 56555 67883
rect 56633 67837 56679 67883
rect 56757 67837 56803 67883
rect 56881 67837 56927 67883
rect 57005 67837 57051 67883
rect 57129 67837 57175 67883
rect 57253 67837 57299 67883
rect 57377 67837 57423 67883
rect 57501 67837 57547 67883
rect 57625 67837 57671 67883
rect 57749 67837 57795 67883
rect 57873 67837 57919 67883
rect 57997 67837 58043 67883
rect 58121 67837 58167 67883
rect 58245 67837 58291 67883
rect 58369 67837 58415 67883
rect 58493 67837 58539 67883
rect 58617 67837 58663 67883
rect 58741 67837 58787 67883
rect 58865 67837 58911 67883
rect 58989 67837 59035 67883
rect 59113 67837 59159 67883
rect 59237 67837 59283 67883
rect 59361 67837 59407 67883
rect 59485 67837 59531 67883
rect 59609 67837 59655 67883
rect 59733 67837 59779 67883
rect 59857 67837 59903 67883
rect 59981 67837 60027 67883
rect 60105 67837 60151 67883
rect 60229 67837 60275 67883
rect 60353 67837 60399 67883
rect 60477 67837 60523 67883
rect 60601 67837 60647 67883
rect 60725 67837 60771 67883
rect 60849 67837 60895 67883
rect 60973 67837 61019 67883
rect 61097 67837 61143 67883
rect 61221 67837 61267 67883
rect 61345 67837 61391 67883
rect 61469 67837 61515 67883
rect 61593 67837 61639 67883
rect 61717 67837 61763 67883
rect 61841 67837 61887 67883
rect 61965 67837 62011 67883
rect 62089 67837 62135 67883
rect 62213 67837 62259 67883
rect 62337 67837 62383 67883
rect 62461 67837 62507 67883
rect 62585 67837 62631 67883
rect 62709 67837 62755 67883
rect 62833 67837 62879 67883
rect 62957 67837 63003 67883
rect 63081 67837 63127 67883
rect 63205 67837 63251 67883
rect 63329 67837 63375 67883
rect 63453 67837 63499 67883
rect 63577 67837 63623 67883
rect 63701 67837 63747 67883
rect 63825 67837 63871 67883
rect 63949 67837 63995 67883
rect 64073 67837 64119 67883
rect 64197 67837 64243 67883
rect 64321 67837 64367 67883
rect 64445 67837 64491 67883
rect 64569 67837 64615 67883
rect 64693 67837 64739 67883
rect 64817 67837 64863 67883
rect 64941 67837 64987 67883
rect 65065 67837 65111 67883
rect 65189 67837 65235 67883
rect 65313 67837 65359 67883
rect 65437 67837 65483 67883
rect 65561 67837 65607 67883
rect 65685 67837 65731 67883
rect 65809 67837 65855 67883
rect 65933 67837 65979 67883
rect 66057 67837 66103 67883
rect 66181 67837 66227 67883
rect 66305 67837 66351 67883
rect 66429 67837 66475 67883
rect 66553 67837 66599 67883
rect 66677 67837 66723 67883
rect 66801 67837 66847 67883
rect 66925 67837 66971 67883
rect 67049 67837 67095 67883
rect 67173 67837 67219 67883
rect 67297 67837 67343 67883
rect 67421 67837 67467 67883
rect 67545 67837 67591 67883
rect 67669 67837 67715 67883
rect 67793 67837 67839 67883
rect 67917 67837 67963 67883
rect 68041 67837 68087 67883
rect 68165 67837 68211 67883
rect 68289 67837 68335 67883
rect 68413 67837 68459 67883
rect 68537 67837 68583 67883
rect 68661 67837 68707 67883
rect 68785 67837 68831 67883
rect 68909 67837 68955 67883
rect 69033 67837 69079 67883
rect 69157 67837 69203 67883
rect 69281 67837 69327 67883
rect 69405 67837 69451 67883
rect 69529 67837 69575 67883
rect 69653 67837 69699 67883
rect 69777 67837 69823 67883
rect 69901 67837 69947 67883
rect 70025 67837 70071 67883
rect 70149 67837 70195 67883
rect 70273 67837 70319 67883
rect 70397 67837 70443 67883
rect 70521 67837 70567 67883
rect 70645 67837 70691 67883
rect 70769 67837 70815 67883
rect 70893 67837 70939 67883
rect 71017 67837 71063 67883
rect 71141 67837 71187 67883
rect 71265 67837 71311 67883
rect 71389 67837 71435 67883
rect 71513 67837 71559 67883
rect 71637 67837 71683 67883
rect 71761 67837 71807 67883
rect 71885 67837 71931 67883
rect 72009 67837 72055 67883
rect 72133 67837 72179 67883
rect 72257 67837 72303 67883
rect 72381 67837 72427 67883
rect 72505 67837 72551 67883
rect 72629 67837 72675 67883
rect 72753 67837 72799 67883
rect 72877 67837 72923 67883
rect 73001 67837 73047 67883
rect 73125 67837 73171 67883
rect 73249 67837 73295 67883
rect 73373 67837 73419 67883
rect 73497 67837 73543 67883
rect 73621 67837 73667 67883
rect 73745 67837 73791 67883
rect 73869 67837 73915 67883
rect 73993 67837 74039 67883
rect 74117 67837 74163 67883
rect 74241 67837 74287 67883
rect 74365 67837 74411 67883
rect 74489 67837 74535 67883
rect 74613 67837 74659 67883
rect 74737 67837 74783 67883
rect 74861 67837 74907 67883
rect 74985 67837 75031 67883
rect 75109 67837 75155 67883
rect 75233 67837 75279 67883
rect 75357 67837 75403 67883
rect 75481 67837 75527 67883
rect 75605 67837 75651 67883
rect 75729 67837 75775 67883
rect 75853 67837 75899 67883
rect 75977 67837 76023 67883
rect 76101 67837 76147 67883
rect 76225 67837 76271 67883
rect 76349 67837 76395 67883
rect 76473 67837 76519 67883
rect 76597 67837 76643 67883
rect 76721 67837 76767 67883
rect 76845 67837 76891 67883
rect 76969 67837 77015 67883
rect 77093 67837 77139 67883
rect 77217 67837 77263 67883
rect 77341 67837 77387 67883
rect 77465 67837 77511 67883
rect 77589 67837 77635 67883
rect 77713 67837 77759 67883
rect 77837 67837 77883 67883
rect 77961 67837 78007 67883
rect 78085 67837 78131 67883
rect 78209 67837 78255 67883
rect 78333 67837 78379 67883
rect 78457 67837 78503 67883
rect 78581 67837 78627 67883
rect 78705 67837 78751 67883
rect 78829 67837 78875 67883
rect 78953 67837 78999 67883
rect 79077 67837 79123 67883
rect 79201 67837 79247 67883
rect 79325 67837 79371 67883
rect 79449 67837 79495 67883
rect 79573 67837 79619 67883
rect 79697 67837 79743 67883
rect 79821 67837 79867 67883
rect 79945 67837 79991 67883
rect 80069 67837 80115 67883
rect 80193 67837 80239 67883
rect 80317 67837 80363 67883
rect 80441 67837 80487 67883
rect 80565 67837 80611 67883
rect 80689 67837 80735 67883
rect 80813 67837 80859 67883
rect 80937 67837 80983 67883
rect 81061 67837 81107 67883
rect 81185 67837 81231 67883
rect 81309 67837 81355 67883
rect 81433 67837 81479 67883
rect 81557 67837 81603 67883
rect 81681 67837 81727 67883
rect 81805 67837 81851 67883
rect 81929 67837 81975 67883
rect 82053 67837 82099 67883
rect 82177 67837 82223 67883
rect 82301 67837 82347 67883
rect 82425 67837 82471 67883
rect 82549 67837 82595 67883
rect 82673 67837 82719 67883
rect 82797 67837 82843 67883
rect 82921 67837 82967 67883
rect 83045 67837 83091 67883
rect 83169 67837 83215 67883
rect 83293 67837 83339 67883
rect 83417 67837 83463 67883
rect 83541 67837 83587 67883
rect 83665 67837 83711 67883
rect 83789 67837 83835 67883
rect 83913 67837 83959 67883
rect 84037 67837 84083 67883
rect 84161 67837 84207 67883
rect 84285 67837 84331 67883
rect 84409 67837 84455 67883
rect 84533 67837 84579 67883
rect 84657 67837 84703 67883
rect 84781 67837 84827 67883
rect 84905 67837 84951 67883
rect 85029 67837 85075 67883
rect 85153 67837 85199 67883
rect 85277 67837 85323 67883
rect 85401 67837 85447 67883
rect 85525 67837 85571 67883
rect 85649 67837 85695 67883
rect 89 67713 135 67759
rect 213 67713 259 67759
rect 337 67713 383 67759
rect 461 67713 507 67759
rect 585 67713 631 67759
rect 709 67713 755 67759
rect 833 67713 879 67759
rect 957 67713 1003 67759
rect 1081 67713 1127 67759
rect 1205 67713 1251 67759
rect 1329 67713 1375 67759
rect 1453 67713 1499 67759
rect 1577 67713 1623 67759
rect 1701 67713 1747 67759
rect 1825 67713 1871 67759
rect 1949 67713 1995 67759
rect 2073 67713 2119 67759
rect 2197 67713 2243 67759
rect 2321 67713 2367 67759
rect 2445 67713 2491 67759
rect 2569 67713 2615 67759
rect 2693 67713 2739 67759
rect 2817 67713 2863 67759
rect 2941 67713 2987 67759
rect 3065 67713 3111 67759
rect 3189 67713 3235 67759
rect 3313 67713 3359 67759
rect 3437 67713 3483 67759
rect 3561 67713 3607 67759
rect 3685 67713 3731 67759
rect 3809 67713 3855 67759
rect 3933 67713 3979 67759
rect 4057 67713 4103 67759
rect 4181 67713 4227 67759
rect 4305 67713 4351 67759
rect 4429 67713 4475 67759
rect 4553 67713 4599 67759
rect 4677 67713 4723 67759
rect 4801 67713 4847 67759
rect 4925 67713 4971 67759
rect 5049 67713 5095 67759
rect 5173 67713 5219 67759
rect 5297 67713 5343 67759
rect 5421 67713 5467 67759
rect 5545 67713 5591 67759
rect 5669 67713 5715 67759
rect 5793 67713 5839 67759
rect 5917 67713 5963 67759
rect 6041 67713 6087 67759
rect 6165 67713 6211 67759
rect 6289 67713 6335 67759
rect 6413 67713 6459 67759
rect 6537 67713 6583 67759
rect 6661 67713 6707 67759
rect 6785 67713 6831 67759
rect 6909 67713 6955 67759
rect 7033 67713 7079 67759
rect 7157 67713 7203 67759
rect 7281 67713 7327 67759
rect 7405 67713 7451 67759
rect 7529 67713 7575 67759
rect 7653 67713 7699 67759
rect 7777 67713 7823 67759
rect 7901 67713 7947 67759
rect 8025 67713 8071 67759
rect 8149 67713 8195 67759
rect 8273 67713 8319 67759
rect 8397 67713 8443 67759
rect 8521 67713 8567 67759
rect 8645 67713 8691 67759
rect 8769 67713 8815 67759
rect 8893 67713 8939 67759
rect 9017 67713 9063 67759
rect 9141 67713 9187 67759
rect 9265 67713 9311 67759
rect 9389 67713 9435 67759
rect 9513 67713 9559 67759
rect 9637 67713 9683 67759
rect 9761 67713 9807 67759
rect 9885 67713 9931 67759
rect 10009 67713 10055 67759
rect 10133 67713 10179 67759
rect 10257 67713 10303 67759
rect 10381 67713 10427 67759
rect 10505 67713 10551 67759
rect 10629 67713 10675 67759
rect 10753 67713 10799 67759
rect 10877 67713 10923 67759
rect 11001 67713 11047 67759
rect 11125 67713 11171 67759
rect 11249 67713 11295 67759
rect 11373 67713 11419 67759
rect 11497 67713 11543 67759
rect 11621 67713 11667 67759
rect 11745 67713 11791 67759
rect 11869 67713 11915 67759
rect 11993 67713 12039 67759
rect 12117 67713 12163 67759
rect 12241 67713 12287 67759
rect 12365 67713 12411 67759
rect 12489 67713 12535 67759
rect 12613 67713 12659 67759
rect 12737 67713 12783 67759
rect 12861 67713 12907 67759
rect 12985 67713 13031 67759
rect 13109 67713 13155 67759
rect 13233 67713 13279 67759
rect 13357 67713 13403 67759
rect 13481 67713 13527 67759
rect 13605 67713 13651 67759
rect 13729 67713 13775 67759
rect 13853 67713 13899 67759
rect 13977 67713 14023 67759
rect 14101 67713 14147 67759
rect 14225 67713 14271 67759
rect 14349 67713 14395 67759
rect 14473 67713 14519 67759
rect 14597 67713 14643 67759
rect 14721 67713 14767 67759
rect 14845 67713 14891 67759
rect 14969 67713 15015 67759
rect 15093 67713 15139 67759
rect 15217 67713 15263 67759
rect 15341 67713 15387 67759
rect 15465 67713 15511 67759
rect 15589 67713 15635 67759
rect 15713 67713 15759 67759
rect 15837 67713 15883 67759
rect 15961 67713 16007 67759
rect 16085 67713 16131 67759
rect 16209 67713 16255 67759
rect 16333 67713 16379 67759
rect 16457 67713 16503 67759
rect 16581 67713 16627 67759
rect 16705 67713 16751 67759
rect 16829 67713 16875 67759
rect 16953 67713 16999 67759
rect 17077 67713 17123 67759
rect 17201 67713 17247 67759
rect 17325 67713 17371 67759
rect 17449 67713 17495 67759
rect 17573 67713 17619 67759
rect 17697 67713 17743 67759
rect 17821 67713 17867 67759
rect 17945 67713 17991 67759
rect 18069 67713 18115 67759
rect 18193 67713 18239 67759
rect 18317 67713 18363 67759
rect 18441 67713 18487 67759
rect 18565 67713 18611 67759
rect 18689 67713 18735 67759
rect 18813 67713 18859 67759
rect 18937 67713 18983 67759
rect 19061 67713 19107 67759
rect 19185 67713 19231 67759
rect 19309 67713 19355 67759
rect 19433 67713 19479 67759
rect 19557 67713 19603 67759
rect 19681 67713 19727 67759
rect 19805 67713 19851 67759
rect 19929 67713 19975 67759
rect 20053 67713 20099 67759
rect 20177 67713 20223 67759
rect 20301 67713 20347 67759
rect 20425 67713 20471 67759
rect 20549 67713 20595 67759
rect 20673 67713 20719 67759
rect 20797 67713 20843 67759
rect 20921 67713 20967 67759
rect 21045 67713 21091 67759
rect 21169 67713 21215 67759
rect 21293 67713 21339 67759
rect 21417 67713 21463 67759
rect 21541 67713 21587 67759
rect 21665 67713 21711 67759
rect 21789 67713 21835 67759
rect 21913 67713 21959 67759
rect 22037 67713 22083 67759
rect 22161 67713 22207 67759
rect 22285 67713 22331 67759
rect 22409 67713 22455 67759
rect 22533 67713 22579 67759
rect 22657 67713 22703 67759
rect 22781 67713 22827 67759
rect 22905 67713 22951 67759
rect 23029 67713 23075 67759
rect 23153 67713 23199 67759
rect 23277 67713 23323 67759
rect 23401 67713 23447 67759
rect 23525 67713 23571 67759
rect 23649 67713 23695 67759
rect 23773 67713 23819 67759
rect 23897 67713 23943 67759
rect 24021 67713 24067 67759
rect 24145 67713 24191 67759
rect 24269 67713 24315 67759
rect 24393 67713 24439 67759
rect 24517 67713 24563 67759
rect 24641 67713 24687 67759
rect 24765 67713 24811 67759
rect 24889 67713 24935 67759
rect 25013 67713 25059 67759
rect 25137 67713 25183 67759
rect 25261 67713 25307 67759
rect 25385 67713 25431 67759
rect 25509 67713 25555 67759
rect 25633 67713 25679 67759
rect 25757 67713 25803 67759
rect 25881 67713 25927 67759
rect 26005 67713 26051 67759
rect 26129 67713 26175 67759
rect 26253 67713 26299 67759
rect 26377 67713 26423 67759
rect 26501 67713 26547 67759
rect 26625 67713 26671 67759
rect 26749 67713 26795 67759
rect 26873 67713 26919 67759
rect 26997 67713 27043 67759
rect 27121 67713 27167 67759
rect 27245 67713 27291 67759
rect 27369 67713 27415 67759
rect 27493 67713 27539 67759
rect 27617 67713 27663 67759
rect 27741 67713 27787 67759
rect 27865 67713 27911 67759
rect 27989 67713 28035 67759
rect 28113 67713 28159 67759
rect 28237 67713 28283 67759
rect 28361 67713 28407 67759
rect 28485 67713 28531 67759
rect 28609 67713 28655 67759
rect 28733 67713 28779 67759
rect 28857 67713 28903 67759
rect 28981 67713 29027 67759
rect 29105 67713 29151 67759
rect 29229 67713 29275 67759
rect 29353 67713 29399 67759
rect 29477 67713 29523 67759
rect 29601 67713 29647 67759
rect 29725 67713 29771 67759
rect 29849 67713 29895 67759
rect 29973 67713 30019 67759
rect 30097 67713 30143 67759
rect 30221 67713 30267 67759
rect 30345 67713 30391 67759
rect 30469 67713 30515 67759
rect 30593 67713 30639 67759
rect 30717 67713 30763 67759
rect 30841 67713 30887 67759
rect 30965 67713 31011 67759
rect 31089 67713 31135 67759
rect 31213 67713 31259 67759
rect 31337 67713 31383 67759
rect 31461 67713 31507 67759
rect 31585 67713 31631 67759
rect 31709 67713 31755 67759
rect 31833 67713 31879 67759
rect 31957 67713 32003 67759
rect 32081 67713 32127 67759
rect 32205 67713 32251 67759
rect 32329 67713 32375 67759
rect 32453 67713 32499 67759
rect 32577 67713 32623 67759
rect 32701 67713 32747 67759
rect 32825 67713 32871 67759
rect 32949 67713 32995 67759
rect 33073 67713 33119 67759
rect 33197 67713 33243 67759
rect 33321 67713 33367 67759
rect 33445 67713 33491 67759
rect 33569 67713 33615 67759
rect 33693 67713 33739 67759
rect 33817 67713 33863 67759
rect 33941 67713 33987 67759
rect 34065 67713 34111 67759
rect 34189 67713 34235 67759
rect 34313 67713 34359 67759
rect 34437 67713 34483 67759
rect 34561 67713 34607 67759
rect 34685 67713 34731 67759
rect 34809 67713 34855 67759
rect 34933 67713 34979 67759
rect 35057 67713 35103 67759
rect 35181 67713 35227 67759
rect 35305 67713 35351 67759
rect 35429 67713 35475 67759
rect 35553 67713 35599 67759
rect 35677 67713 35723 67759
rect 35801 67713 35847 67759
rect 35925 67713 35971 67759
rect 36049 67713 36095 67759
rect 36173 67713 36219 67759
rect 36297 67713 36343 67759
rect 36421 67713 36467 67759
rect 36545 67713 36591 67759
rect 36669 67713 36715 67759
rect 36793 67713 36839 67759
rect 36917 67713 36963 67759
rect 37041 67713 37087 67759
rect 37165 67713 37211 67759
rect 37289 67713 37335 67759
rect 37413 67713 37459 67759
rect 37537 67713 37583 67759
rect 37661 67713 37707 67759
rect 37785 67713 37831 67759
rect 37909 67713 37955 67759
rect 38033 67713 38079 67759
rect 38157 67713 38203 67759
rect 38281 67713 38327 67759
rect 38405 67713 38451 67759
rect 38529 67713 38575 67759
rect 38653 67713 38699 67759
rect 38777 67713 38823 67759
rect 38901 67713 38947 67759
rect 39025 67713 39071 67759
rect 39149 67713 39195 67759
rect 39273 67713 39319 67759
rect 39397 67713 39443 67759
rect 39521 67713 39567 67759
rect 39645 67713 39691 67759
rect 39769 67713 39815 67759
rect 39893 67713 39939 67759
rect 40017 67713 40063 67759
rect 40141 67713 40187 67759
rect 40265 67713 40311 67759
rect 40389 67713 40435 67759
rect 40513 67713 40559 67759
rect 40637 67713 40683 67759
rect 40761 67713 40807 67759
rect 40885 67713 40931 67759
rect 41009 67713 41055 67759
rect 41133 67713 41179 67759
rect 41257 67713 41303 67759
rect 41381 67713 41427 67759
rect 41505 67713 41551 67759
rect 41629 67713 41675 67759
rect 41753 67713 41799 67759
rect 41877 67713 41923 67759
rect 42001 67713 42047 67759
rect 42125 67713 42171 67759
rect 42249 67713 42295 67759
rect 42373 67713 42419 67759
rect 42497 67713 42543 67759
rect 42621 67713 42667 67759
rect 42745 67713 42791 67759
rect 42869 67713 42915 67759
rect 42993 67713 43039 67759
rect 43117 67713 43163 67759
rect 43241 67713 43287 67759
rect 43365 67713 43411 67759
rect 43489 67713 43535 67759
rect 43613 67713 43659 67759
rect 43737 67713 43783 67759
rect 43861 67713 43907 67759
rect 43985 67713 44031 67759
rect 44109 67713 44155 67759
rect 44233 67713 44279 67759
rect 44357 67713 44403 67759
rect 44481 67713 44527 67759
rect 44605 67713 44651 67759
rect 44729 67713 44775 67759
rect 44853 67713 44899 67759
rect 44977 67713 45023 67759
rect 45101 67713 45147 67759
rect 45225 67713 45271 67759
rect 45349 67713 45395 67759
rect 45473 67713 45519 67759
rect 45597 67713 45643 67759
rect 45721 67713 45767 67759
rect 45845 67713 45891 67759
rect 45969 67713 46015 67759
rect 46093 67713 46139 67759
rect 46217 67713 46263 67759
rect 46341 67713 46387 67759
rect 46465 67713 46511 67759
rect 46589 67713 46635 67759
rect 46713 67713 46759 67759
rect 46837 67713 46883 67759
rect 46961 67713 47007 67759
rect 47085 67713 47131 67759
rect 47209 67713 47255 67759
rect 47333 67713 47379 67759
rect 47457 67713 47503 67759
rect 47581 67713 47627 67759
rect 47705 67713 47751 67759
rect 47829 67713 47875 67759
rect 47953 67713 47999 67759
rect 48077 67713 48123 67759
rect 48201 67713 48247 67759
rect 48325 67713 48371 67759
rect 48449 67713 48495 67759
rect 48573 67713 48619 67759
rect 48697 67713 48743 67759
rect 48821 67713 48867 67759
rect 48945 67713 48991 67759
rect 49069 67713 49115 67759
rect 49193 67713 49239 67759
rect 49317 67713 49363 67759
rect 49441 67713 49487 67759
rect 49565 67713 49611 67759
rect 49689 67713 49735 67759
rect 49813 67713 49859 67759
rect 49937 67713 49983 67759
rect 50061 67713 50107 67759
rect 50185 67713 50231 67759
rect 50309 67713 50355 67759
rect 50433 67713 50479 67759
rect 50557 67713 50603 67759
rect 50681 67713 50727 67759
rect 50805 67713 50851 67759
rect 50929 67713 50975 67759
rect 51053 67713 51099 67759
rect 51177 67713 51223 67759
rect 51301 67713 51347 67759
rect 51425 67713 51471 67759
rect 51549 67713 51595 67759
rect 51673 67713 51719 67759
rect 51797 67713 51843 67759
rect 51921 67713 51967 67759
rect 52045 67713 52091 67759
rect 52169 67713 52215 67759
rect 52293 67713 52339 67759
rect 52417 67713 52463 67759
rect 52541 67713 52587 67759
rect 52665 67713 52711 67759
rect 52789 67713 52835 67759
rect 52913 67713 52959 67759
rect 53037 67713 53083 67759
rect 53161 67713 53207 67759
rect 53285 67713 53331 67759
rect 53409 67713 53455 67759
rect 53533 67713 53579 67759
rect 53657 67713 53703 67759
rect 53781 67713 53827 67759
rect 53905 67713 53951 67759
rect 54029 67713 54075 67759
rect 54153 67713 54199 67759
rect 54277 67713 54323 67759
rect 54401 67713 54447 67759
rect 54525 67713 54571 67759
rect 54649 67713 54695 67759
rect 54773 67713 54819 67759
rect 54897 67713 54943 67759
rect 55021 67713 55067 67759
rect 55145 67713 55191 67759
rect 55269 67713 55315 67759
rect 55393 67713 55439 67759
rect 55517 67713 55563 67759
rect 55641 67713 55687 67759
rect 55765 67713 55811 67759
rect 55889 67713 55935 67759
rect 56013 67713 56059 67759
rect 56137 67713 56183 67759
rect 56261 67713 56307 67759
rect 56385 67713 56431 67759
rect 56509 67713 56555 67759
rect 56633 67713 56679 67759
rect 56757 67713 56803 67759
rect 56881 67713 56927 67759
rect 57005 67713 57051 67759
rect 57129 67713 57175 67759
rect 57253 67713 57299 67759
rect 57377 67713 57423 67759
rect 57501 67713 57547 67759
rect 57625 67713 57671 67759
rect 57749 67713 57795 67759
rect 57873 67713 57919 67759
rect 57997 67713 58043 67759
rect 58121 67713 58167 67759
rect 58245 67713 58291 67759
rect 58369 67713 58415 67759
rect 58493 67713 58539 67759
rect 58617 67713 58663 67759
rect 58741 67713 58787 67759
rect 58865 67713 58911 67759
rect 58989 67713 59035 67759
rect 59113 67713 59159 67759
rect 59237 67713 59283 67759
rect 59361 67713 59407 67759
rect 59485 67713 59531 67759
rect 59609 67713 59655 67759
rect 59733 67713 59779 67759
rect 59857 67713 59903 67759
rect 59981 67713 60027 67759
rect 60105 67713 60151 67759
rect 60229 67713 60275 67759
rect 60353 67713 60399 67759
rect 60477 67713 60523 67759
rect 60601 67713 60647 67759
rect 60725 67713 60771 67759
rect 60849 67713 60895 67759
rect 60973 67713 61019 67759
rect 61097 67713 61143 67759
rect 61221 67713 61267 67759
rect 61345 67713 61391 67759
rect 61469 67713 61515 67759
rect 61593 67713 61639 67759
rect 61717 67713 61763 67759
rect 61841 67713 61887 67759
rect 61965 67713 62011 67759
rect 62089 67713 62135 67759
rect 62213 67713 62259 67759
rect 62337 67713 62383 67759
rect 62461 67713 62507 67759
rect 62585 67713 62631 67759
rect 62709 67713 62755 67759
rect 62833 67713 62879 67759
rect 62957 67713 63003 67759
rect 63081 67713 63127 67759
rect 63205 67713 63251 67759
rect 63329 67713 63375 67759
rect 63453 67713 63499 67759
rect 63577 67713 63623 67759
rect 63701 67713 63747 67759
rect 63825 67713 63871 67759
rect 63949 67713 63995 67759
rect 64073 67713 64119 67759
rect 64197 67713 64243 67759
rect 64321 67713 64367 67759
rect 64445 67713 64491 67759
rect 64569 67713 64615 67759
rect 64693 67713 64739 67759
rect 64817 67713 64863 67759
rect 64941 67713 64987 67759
rect 65065 67713 65111 67759
rect 65189 67713 65235 67759
rect 65313 67713 65359 67759
rect 65437 67713 65483 67759
rect 65561 67713 65607 67759
rect 65685 67713 65731 67759
rect 65809 67713 65855 67759
rect 65933 67713 65979 67759
rect 66057 67713 66103 67759
rect 66181 67713 66227 67759
rect 66305 67713 66351 67759
rect 66429 67713 66475 67759
rect 66553 67713 66599 67759
rect 66677 67713 66723 67759
rect 66801 67713 66847 67759
rect 66925 67713 66971 67759
rect 67049 67713 67095 67759
rect 67173 67713 67219 67759
rect 67297 67713 67343 67759
rect 67421 67713 67467 67759
rect 67545 67713 67591 67759
rect 67669 67713 67715 67759
rect 67793 67713 67839 67759
rect 67917 67713 67963 67759
rect 68041 67713 68087 67759
rect 68165 67713 68211 67759
rect 68289 67713 68335 67759
rect 68413 67713 68459 67759
rect 68537 67713 68583 67759
rect 68661 67713 68707 67759
rect 68785 67713 68831 67759
rect 68909 67713 68955 67759
rect 69033 67713 69079 67759
rect 69157 67713 69203 67759
rect 69281 67713 69327 67759
rect 69405 67713 69451 67759
rect 69529 67713 69575 67759
rect 69653 67713 69699 67759
rect 69777 67713 69823 67759
rect 69901 67713 69947 67759
rect 70025 67713 70071 67759
rect 70149 67713 70195 67759
rect 70273 67713 70319 67759
rect 70397 67713 70443 67759
rect 70521 67713 70567 67759
rect 70645 67713 70691 67759
rect 70769 67713 70815 67759
rect 70893 67713 70939 67759
rect 71017 67713 71063 67759
rect 71141 67713 71187 67759
rect 71265 67713 71311 67759
rect 71389 67713 71435 67759
rect 71513 67713 71559 67759
rect 71637 67713 71683 67759
rect 71761 67713 71807 67759
rect 71885 67713 71931 67759
rect 72009 67713 72055 67759
rect 72133 67713 72179 67759
rect 72257 67713 72303 67759
rect 72381 67713 72427 67759
rect 72505 67713 72551 67759
rect 72629 67713 72675 67759
rect 72753 67713 72799 67759
rect 72877 67713 72923 67759
rect 73001 67713 73047 67759
rect 73125 67713 73171 67759
rect 73249 67713 73295 67759
rect 73373 67713 73419 67759
rect 73497 67713 73543 67759
rect 73621 67713 73667 67759
rect 73745 67713 73791 67759
rect 73869 67713 73915 67759
rect 73993 67713 74039 67759
rect 74117 67713 74163 67759
rect 74241 67713 74287 67759
rect 74365 67713 74411 67759
rect 74489 67713 74535 67759
rect 74613 67713 74659 67759
rect 74737 67713 74783 67759
rect 74861 67713 74907 67759
rect 74985 67713 75031 67759
rect 75109 67713 75155 67759
rect 75233 67713 75279 67759
rect 75357 67713 75403 67759
rect 75481 67713 75527 67759
rect 75605 67713 75651 67759
rect 75729 67713 75775 67759
rect 75853 67713 75899 67759
rect 75977 67713 76023 67759
rect 76101 67713 76147 67759
rect 76225 67713 76271 67759
rect 76349 67713 76395 67759
rect 76473 67713 76519 67759
rect 76597 67713 76643 67759
rect 76721 67713 76767 67759
rect 76845 67713 76891 67759
rect 76969 67713 77015 67759
rect 77093 67713 77139 67759
rect 77217 67713 77263 67759
rect 77341 67713 77387 67759
rect 77465 67713 77511 67759
rect 77589 67713 77635 67759
rect 77713 67713 77759 67759
rect 77837 67713 77883 67759
rect 77961 67713 78007 67759
rect 78085 67713 78131 67759
rect 78209 67713 78255 67759
rect 78333 67713 78379 67759
rect 78457 67713 78503 67759
rect 78581 67713 78627 67759
rect 78705 67713 78751 67759
rect 78829 67713 78875 67759
rect 78953 67713 78999 67759
rect 79077 67713 79123 67759
rect 79201 67713 79247 67759
rect 79325 67713 79371 67759
rect 79449 67713 79495 67759
rect 79573 67713 79619 67759
rect 79697 67713 79743 67759
rect 79821 67713 79867 67759
rect 79945 67713 79991 67759
rect 80069 67713 80115 67759
rect 80193 67713 80239 67759
rect 80317 67713 80363 67759
rect 80441 67713 80487 67759
rect 80565 67713 80611 67759
rect 80689 67713 80735 67759
rect 80813 67713 80859 67759
rect 80937 67713 80983 67759
rect 81061 67713 81107 67759
rect 81185 67713 81231 67759
rect 81309 67713 81355 67759
rect 81433 67713 81479 67759
rect 81557 67713 81603 67759
rect 81681 67713 81727 67759
rect 81805 67713 81851 67759
rect 81929 67713 81975 67759
rect 82053 67713 82099 67759
rect 82177 67713 82223 67759
rect 82301 67713 82347 67759
rect 82425 67713 82471 67759
rect 82549 67713 82595 67759
rect 82673 67713 82719 67759
rect 82797 67713 82843 67759
rect 82921 67713 82967 67759
rect 83045 67713 83091 67759
rect 83169 67713 83215 67759
rect 83293 67713 83339 67759
rect 83417 67713 83463 67759
rect 83541 67713 83587 67759
rect 83665 67713 83711 67759
rect 83789 67713 83835 67759
rect 83913 67713 83959 67759
rect 84037 67713 84083 67759
rect 84161 67713 84207 67759
rect 84285 67713 84331 67759
rect 84409 67713 84455 67759
rect 84533 67713 84579 67759
rect 84657 67713 84703 67759
rect 84781 67713 84827 67759
rect 84905 67713 84951 67759
rect 85029 67713 85075 67759
rect 85153 67713 85199 67759
rect 85277 67713 85323 67759
rect 85401 67713 85447 67759
rect 85525 67713 85571 67759
rect 85649 67713 85695 67759
rect 89 67589 135 67635
rect 213 67589 259 67635
rect 337 67589 383 67635
rect 461 67589 507 67635
rect 585 67589 631 67635
rect 709 67589 755 67635
rect 833 67589 879 67635
rect 957 67589 1003 67635
rect 1081 67589 1127 67635
rect 1205 67589 1251 67635
rect 1329 67589 1375 67635
rect 1453 67589 1499 67635
rect 1577 67589 1623 67635
rect 1701 67589 1747 67635
rect 1825 67589 1871 67635
rect 1949 67589 1995 67635
rect 2073 67589 2119 67635
rect 2197 67589 2243 67635
rect 2321 67589 2367 67635
rect 2445 67589 2491 67635
rect 2569 67589 2615 67635
rect 2693 67589 2739 67635
rect 2817 67589 2863 67635
rect 2941 67589 2987 67635
rect 3065 67589 3111 67635
rect 3189 67589 3235 67635
rect 3313 67589 3359 67635
rect 3437 67589 3483 67635
rect 3561 67589 3607 67635
rect 3685 67589 3731 67635
rect 3809 67589 3855 67635
rect 3933 67589 3979 67635
rect 4057 67589 4103 67635
rect 4181 67589 4227 67635
rect 4305 67589 4351 67635
rect 4429 67589 4475 67635
rect 4553 67589 4599 67635
rect 4677 67589 4723 67635
rect 4801 67589 4847 67635
rect 4925 67589 4971 67635
rect 5049 67589 5095 67635
rect 5173 67589 5219 67635
rect 5297 67589 5343 67635
rect 5421 67589 5467 67635
rect 5545 67589 5591 67635
rect 5669 67589 5715 67635
rect 5793 67589 5839 67635
rect 5917 67589 5963 67635
rect 6041 67589 6087 67635
rect 6165 67589 6211 67635
rect 6289 67589 6335 67635
rect 6413 67589 6459 67635
rect 6537 67589 6583 67635
rect 6661 67589 6707 67635
rect 6785 67589 6831 67635
rect 6909 67589 6955 67635
rect 7033 67589 7079 67635
rect 7157 67589 7203 67635
rect 7281 67589 7327 67635
rect 7405 67589 7451 67635
rect 7529 67589 7575 67635
rect 7653 67589 7699 67635
rect 7777 67589 7823 67635
rect 7901 67589 7947 67635
rect 8025 67589 8071 67635
rect 8149 67589 8195 67635
rect 8273 67589 8319 67635
rect 8397 67589 8443 67635
rect 8521 67589 8567 67635
rect 8645 67589 8691 67635
rect 8769 67589 8815 67635
rect 8893 67589 8939 67635
rect 9017 67589 9063 67635
rect 9141 67589 9187 67635
rect 9265 67589 9311 67635
rect 9389 67589 9435 67635
rect 9513 67589 9559 67635
rect 9637 67589 9683 67635
rect 9761 67589 9807 67635
rect 9885 67589 9931 67635
rect 10009 67589 10055 67635
rect 10133 67589 10179 67635
rect 10257 67589 10303 67635
rect 10381 67589 10427 67635
rect 10505 67589 10551 67635
rect 10629 67589 10675 67635
rect 10753 67589 10799 67635
rect 10877 67589 10923 67635
rect 11001 67589 11047 67635
rect 11125 67589 11171 67635
rect 11249 67589 11295 67635
rect 11373 67589 11419 67635
rect 11497 67589 11543 67635
rect 11621 67589 11667 67635
rect 11745 67589 11791 67635
rect 11869 67589 11915 67635
rect 11993 67589 12039 67635
rect 12117 67589 12163 67635
rect 12241 67589 12287 67635
rect 12365 67589 12411 67635
rect 12489 67589 12535 67635
rect 12613 67589 12659 67635
rect 12737 67589 12783 67635
rect 12861 67589 12907 67635
rect 12985 67589 13031 67635
rect 13109 67589 13155 67635
rect 13233 67589 13279 67635
rect 13357 67589 13403 67635
rect 13481 67589 13527 67635
rect 13605 67589 13651 67635
rect 13729 67589 13775 67635
rect 13853 67589 13899 67635
rect 13977 67589 14023 67635
rect 14101 67589 14147 67635
rect 14225 67589 14271 67635
rect 14349 67589 14395 67635
rect 14473 67589 14519 67635
rect 14597 67589 14643 67635
rect 14721 67589 14767 67635
rect 14845 67589 14891 67635
rect 14969 67589 15015 67635
rect 15093 67589 15139 67635
rect 15217 67589 15263 67635
rect 15341 67589 15387 67635
rect 15465 67589 15511 67635
rect 15589 67589 15635 67635
rect 15713 67589 15759 67635
rect 15837 67589 15883 67635
rect 15961 67589 16007 67635
rect 16085 67589 16131 67635
rect 16209 67589 16255 67635
rect 16333 67589 16379 67635
rect 16457 67589 16503 67635
rect 16581 67589 16627 67635
rect 16705 67589 16751 67635
rect 16829 67589 16875 67635
rect 16953 67589 16999 67635
rect 17077 67589 17123 67635
rect 17201 67589 17247 67635
rect 17325 67589 17371 67635
rect 17449 67589 17495 67635
rect 17573 67589 17619 67635
rect 17697 67589 17743 67635
rect 17821 67589 17867 67635
rect 17945 67589 17991 67635
rect 18069 67589 18115 67635
rect 18193 67589 18239 67635
rect 18317 67589 18363 67635
rect 18441 67589 18487 67635
rect 18565 67589 18611 67635
rect 18689 67589 18735 67635
rect 18813 67589 18859 67635
rect 18937 67589 18983 67635
rect 19061 67589 19107 67635
rect 19185 67589 19231 67635
rect 19309 67589 19355 67635
rect 19433 67589 19479 67635
rect 19557 67589 19603 67635
rect 19681 67589 19727 67635
rect 19805 67589 19851 67635
rect 19929 67589 19975 67635
rect 20053 67589 20099 67635
rect 20177 67589 20223 67635
rect 20301 67589 20347 67635
rect 20425 67589 20471 67635
rect 20549 67589 20595 67635
rect 20673 67589 20719 67635
rect 20797 67589 20843 67635
rect 20921 67589 20967 67635
rect 21045 67589 21091 67635
rect 21169 67589 21215 67635
rect 21293 67589 21339 67635
rect 21417 67589 21463 67635
rect 21541 67589 21587 67635
rect 21665 67589 21711 67635
rect 21789 67589 21835 67635
rect 21913 67589 21959 67635
rect 22037 67589 22083 67635
rect 22161 67589 22207 67635
rect 22285 67589 22331 67635
rect 22409 67589 22455 67635
rect 22533 67589 22579 67635
rect 22657 67589 22703 67635
rect 22781 67589 22827 67635
rect 22905 67589 22951 67635
rect 23029 67589 23075 67635
rect 23153 67589 23199 67635
rect 23277 67589 23323 67635
rect 23401 67589 23447 67635
rect 23525 67589 23571 67635
rect 23649 67589 23695 67635
rect 23773 67589 23819 67635
rect 23897 67589 23943 67635
rect 24021 67589 24067 67635
rect 24145 67589 24191 67635
rect 24269 67589 24315 67635
rect 24393 67589 24439 67635
rect 24517 67589 24563 67635
rect 24641 67589 24687 67635
rect 24765 67589 24811 67635
rect 24889 67589 24935 67635
rect 25013 67589 25059 67635
rect 25137 67589 25183 67635
rect 25261 67589 25307 67635
rect 25385 67589 25431 67635
rect 25509 67589 25555 67635
rect 25633 67589 25679 67635
rect 25757 67589 25803 67635
rect 25881 67589 25927 67635
rect 26005 67589 26051 67635
rect 26129 67589 26175 67635
rect 26253 67589 26299 67635
rect 26377 67589 26423 67635
rect 26501 67589 26547 67635
rect 26625 67589 26671 67635
rect 26749 67589 26795 67635
rect 26873 67589 26919 67635
rect 26997 67589 27043 67635
rect 27121 67589 27167 67635
rect 27245 67589 27291 67635
rect 27369 67589 27415 67635
rect 27493 67589 27539 67635
rect 27617 67589 27663 67635
rect 27741 67589 27787 67635
rect 27865 67589 27911 67635
rect 27989 67589 28035 67635
rect 28113 67589 28159 67635
rect 28237 67589 28283 67635
rect 28361 67589 28407 67635
rect 28485 67589 28531 67635
rect 28609 67589 28655 67635
rect 28733 67589 28779 67635
rect 28857 67589 28903 67635
rect 28981 67589 29027 67635
rect 29105 67589 29151 67635
rect 29229 67589 29275 67635
rect 29353 67589 29399 67635
rect 29477 67589 29523 67635
rect 29601 67589 29647 67635
rect 29725 67589 29771 67635
rect 29849 67589 29895 67635
rect 29973 67589 30019 67635
rect 30097 67589 30143 67635
rect 30221 67589 30267 67635
rect 30345 67589 30391 67635
rect 30469 67589 30515 67635
rect 30593 67589 30639 67635
rect 30717 67589 30763 67635
rect 30841 67589 30887 67635
rect 30965 67589 31011 67635
rect 31089 67589 31135 67635
rect 31213 67589 31259 67635
rect 31337 67589 31383 67635
rect 31461 67589 31507 67635
rect 31585 67589 31631 67635
rect 31709 67589 31755 67635
rect 31833 67589 31879 67635
rect 31957 67589 32003 67635
rect 32081 67589 32127 67635
rect 32205 67589 32251 67635
rect 32329 67589 32375 67635
rect 32453 67589 32499 67635
rect 32577 67589 32623 67635
rect 32701 67589 32747 67635
rect 32825 67589 32871 67635
rect 32949 67589 32995 67635
rect 33073 67589 33119 67635
rect 33197 67589 33243 67635
rect 33321 67589 33367 67635
rect 33445 67589 33491 67635
rect 33569 67589 33615 67635
rect 33693 67589 33739 67635
rect 33817 67589 33863 67635
rect 33941 67589 33987 67635
rect 34065 67589 34111 67635
rect 34189 67589 34235 67635
rect 34313 67589 34359 67635
rect 34437 67589 34483 67635
rect 34561 67589 34607 67635
rect 34685 67589 34731 67635
rect 34809 67589 34855 67635
rect 34933 67589 34979 67635
rect 35057 67589 35103 67635
rect 35181 67589 35227 67635
rect 35305 67589 35351 67635
rect 35429 67589 35475 67635
rect 35553 67589 35599 67635
rect 35677 67589 35723 67635
rect 35801 67589 35847 67635
rect 35925 67589 35971 67635
rect 36049 67589 36095 67635
rect 36173 67589 36219 67635
rect 36297 67589 36343 67635
rect 36421 67589 36467 67635
rect 36545 67589 36591 67635
rect 36669 67589 36715 67635
rect 36793 67589 36839 67635
rect 36917 67589 36963 67635
rect 37041 67589 37087 67635
rect 37165 67589 37211 67635
rect 37289 67589 37335 67635
rect 37413 67589 37459 67635
rect 37537 67589 37583 67635
rect 37661 67589 37707 67635
rect 37785 67589 37831 67635
rect 37909 67589 37955 67635
rect 38033 67589 38079 67635
rect 38157 67589 38203 67635
rect 38281 67589 38327 67635
rect 38405 67589 38451 67635
rect 38529 67589 38575 67635
rect 38653 67589 38699 67635
rect 38777 67589 38823 67635
rect 38901 67589 38947 67635
rect 39025 67589 39071 67635
rect 39149 67589 39195 67635
rect 39273 67589 39319 67635
rect 39397 67589 39443 67635
rect 39521 67589 39567 67635
rect 39645 67589 39691 67635
rect 39769 67589 39815 67635
rect 39893 67589 39939 67635
rect 40017 67589 40063 67635
rect 40141 67589 40187 67635
rect 40265 67589 40311 67635
rect 40389 67589 40435 67635
rect 40513 67589 40559 67635
rect 40637 67589 40683 67635
rect 40761 67589 40807 67635
rect 40885 67589 40931 67635
rect 41009 67589 41055 67635
rect 41133 67589 41179 67635
rect 41257 67589 41303 67635
rect 41381 67589 41427 67635
rect 41505 67589 41551 67635
rect 41629 67589 41675 67635
rect 41753 67589 41799 67635
rect 41877 67589 41923 67635
rect 42001 67589 42047 67635
rect 42125 67589 42171 67635
rect 42249 67589 42295 67635
rect 42373 67589 42419 67635
rect 42497 67589 42543 67635
rect 42621 67589 42667 67635
rect 42745 67589 42791 67635
rect 42869 67589 42915 67635
rect 42993 67589 43039 67635
rect 43117 67589 43163 67635
rect 43241 67589 43287 67635
rect 43365 67589 43411 67635
rect 43489 67589 43535 67635
rect 43613 67589 43659 67635
rect 43737 67589 43783 67635
rect 43861 67589 43907 67635
rect 43985 67589 44031 67635
rect 44109 67589 44155 67635
rect 44233 67589 44279 67635
rect 44357 67589 44403 67635
rect 44481 67589 44527 67635
rect 44605 67589 44651 67635
rect 44729 67589 44775 67635
rect 44853 67589 44899 67635
rect 44977 67589 45023 67635
rect 45101 67589 45147 67635
rect 45225 67589 45271 67635
rect 45349 67589 45395 67635
rect 45473 67589 45519 67635
rect 45597 67589 45643 67635
rect 45721 67589 45767 67635
rect 45845 67589 45891 67635
rect 45969 67589 46015 67635
rect 46093 67589 46139 67635
rect 46217 67589 46263 67635
rect 46341 67589 46387 67635
rect 46465 67589 46511 67635
rect 46589 67589 46635 67635
rect 46713 67589 46759 67635
rect 46837 67589 46883 67635
rect 46961 67589 47007 67635
rect 47085 67589 47131 67635
rect 47209 67589 47255 67635
rect 47333 67589 47379 67635
rect 47457 67589 47503 67635
rect 47581 67589 47627 67635
rect 47705 67589 47751 67635
rect 47829 67589 47875 67635
rect 47953 67589 47999 67635
rect 48077 67589 48123 67635
rect 48201 67589 48247 67635
rect 48325 67589 48371 67635
rect 48449 67589 48495 67635
rect 48573 67589 48619 67635
rect 48697 67589 48743 67635
rect 48821 67589 48867 67635
rect 48945 67589 48991 67635
rect 49069 67589 49115 67635
rect 49193 67589 49239 67635
rect 49317 67589 49363 67635
rect 49441 67589 49487 67635
rect 49565 67589 49611 67635
rect 49689 67589 49735 67635
rect 49813 67589 49859 67635
rect 49937 67589 49983 67635
rect 50061 67589 50107 67635
rect 50185 67589 50231 67635
rect 50309 67589 50355 67635
rect 50433 67589 50479 67635
rect 50557 67589 50603 67635
rect 50681 67589 50727 67635
rect 50805 67589 50851 67635
rect 50929 67589 50975 67635
rect 51053 67589 51099 67635
rect 51177 67589 51223 67635
rect 51301 67589 51347 67635
rect 51425 67589 51471 67635
rect 51549 67589 51595 67635
rect 51673 67589 51719 67635
rect 51797 67589 51843 67635
rect 51921 67589 51967 67635
rect 52045 67589 52091 67635
rect 52169 67589 52215 67635
rect 52293 67589 52339 67635
rect 52417 67589 52463 67635
rect 52541 67589 52587 67635
rect 52665 67589 52711 67635
rect 52789 67589 52835 67635
rect 52913 67589 52959 67635
rect 53037 67589 53083 67635
rect 53161 67589 53207 67635
rect 53285 67589 53331 67635
rect 53409 67589 53455 67635
rect 53533 67589 53579 67635
rect 53657 67589 53703 67635
rect 53781 67589 53827 67635
rect 53905 67589 53951 67635
rect 54029 67589 54075 67635
rect 54153 67589 54199 67635
rect 54277 67589 54323 67635
rect 54401 67589 54447 67635
rect 54525 67589 54571 67635
rect 54649 67589 54695 67635
rect 54773 67589 54819 67635
rect 54897 67589 54943 67635
rect 55021 67589 55067 67635
rect 55145 67589 55191 67635
rect 55269 67589 55315 67635
rect 55393 67589 55439 67635
rect 55517 67589 55563 67635
rect 55641 67589 55687 67635
rect 55765 67589 55811 67635
rect 55889 67589 55935 67635
rect 56013 67589 56059 67635
rect 56137 67589 56183 67635
rect 56261 67589 56307 67635
rect 56385 67589 56431 67635
rect 56509 67589 56555 67635
rect 56633 67589 56679 67635
rect 56757 67589 56803 67635
rect 56881 67589 56927 67635
rect 57005 67589 57051 67635
rect 57129 67589 57175 67635
rect 57253 67589 57299 67635
rect 57377 67589 57423 67635
rect 57501 67589 57547 67635
rect 57625 67589 57671 67635
rect 57749 67589 57795 67635
rect 57873 67589 57919 67635
rect 57997 67589 58043 67635
rect 58121 67589 58167 67635
rect 58245 67589 58291 67635
rect 58369 67589 58415 67635
rect 58493 67589 58539 67635
rect 58617 67589 58663 67635
rect 58741 67589 58787 67635
rect 58865 67589 58911 67635
rect 58989 67589 59035 67635
rect 59113 67589 59159 67635
rect 59237 67589 59283 67635
rect 59361 67589 59407 67635
rect 59485 67589 59531 67635
rect 59609 67589 59655 67635
rect 59733 67589 59779 67635
rect 59857 67589 59903 67635
rect 59981 67589 60027 67635
rect 60105 67589 60151 67635
rect 60229 67589 60275 67635
rect 60353 67589 60399 67635
rect 60477 67589 60523 67635
rect 60601 67589 60647 67635
rect 60725 67589 60771 67635
rect 60849 67589 60895 67635
rect 60973 67589 61019 67635
rect 61097 67589 61143 67635
rect 61221 67589 61267 67635
rect 61345 67589 61391 67635
rect 61469 67589 61515 67635
rect 61593 67589 61639 67635
rect 61717 67589 61763 67635
rect 61841 67589 61887 67635
rect 61965 67589 62011 67635
rect 62089 67589 62135 67635
rect 62213 67589 62259 67635
rect 62337 67589 62383 67635
rect 62461 67589 62507 67635
rect 62585 67589 62631 67635
rect 62709 67589 62755 67635
rect 62833 67589 62879 67635
rect 62957 67589 63003 67635
rect 63081 67589 63127 67635
rect 63205 67589 63251 67635
rect 63329 67589 63375 67635
rect 63453 67589 63499 67635
rect 63577 67589 63623 67635
rect 63701 67589 63747 67635
rect 63825 67589 63871 67635
rect 63949 67589 63995 67635
rect 64073 67589 64119 67635
rect 64197 67589 64243 67635
rect 64321 67589 64367 67635
rect 64445 67589 64491 67635
rect 64569 67589 64615 67635
rect 64693 67589 64739 67635
rect 64817 67589 64863 67635
rect 64941 67589 64987 67635
rect 65065 67589 65111 67635
rect 65189 67589 65235 67635
rect 65313 67589 65359 67635
rect 65437 67589 65483 67635
rect 65561 67589 65607 67635
rect 65685 67589 65731 67635
rect 65809 67589 65855 67635
rect 65933 67589 65979 67635
rect 66057 67589 66103 67635
rect 66181 67589 66227 67635
rect 66305 67589 66351 67635
rect 66429 67589 66475 67635
rect 66553 67589 66599 67635
rect 66677 67589 66723 67635
rect 66801 67589 66847 67635
rect 66925 67589 66971 67635
rect 67049 67589 67095 67635
rect 67173 67589 67219 67635
rect 67297 67589 67343 67635
rect 67421 67589 67467 67635
rect 67545 67589 67591 67635
rect 67669 67589 67715 67635
rect 67793 67589 67839 67635
rect 67917 67589 67963 67635
rect 68041 67589 68087 67635
rect 68165 67589 68211 67635
rect 68289 67589 68335 67635
rect 68413 67589 68459 67635
rect 68537 67589 68583 67635
rect 68661 67589 68707 67635
rect 68785 67589 68831 67635
rect 68909 67589 68955 67635
rect 69033 67589 69079 67635
rect 69157 67589 69203 67635
rect 69281 67589 69327 67635
rect 69405 67589 69451 67635
rect 69529 67589 69575 67635
rect 69653 67589 69699 67635
rect 69777 67589 69823 67635
rect 69901 67589 69947 67635
rect 70025 67589 70071 67635
rect 70149 67589 70195 67635
rect 70273 67589 70319 67635
rect 70397 67589 70443 67635
rect 70521 67589 70567 67635
rect 70645 67589 70691 67635
rect 70769 67589 70815 67635
rect 70893 67589 70939 67635
rect 71017 67589 71063 67635
rect 71141 67589 71187 67635
rect 71265 67589 71311 67635
rect 71389 67589 71435 67635
rect 71513 67589 71559 67635
rect 71637 67589 71683 67635
rect 71761 67589 71807 67635
rect 71885 67589 71931 67635
rect 72009 67589 72055 67635
rect 72133 67589 72179 67635
rect 72257 67589 72303 67635
rect 72381 67589 72427 67635
rect 72505 67589 72551 67635
rect 72629 67589 72675 67635
rect 72753 67589 72799 67635
rect 72877 67589 72923 67635
rect 73001 67589 73047 67635
rect 73125 67589 73171 67635
rect 73249 67589 73295 67635
rect 73373 67589 73419 67635
rect 73497 67589 73543 67635
rect 73621 67589 73667 67635
rect 73745 67589 73791 67635
rect 73869 67589 73915 67635
rect 73993 67589 74039 67635
rect 74117 67589 74163 67635
rect 74241 67589 74287 67635
rect 74365 67589 74411 67635
rect 74489 67589 74535 67635
rect 74613 67589 74659 67635
rect 74737 67589 74783 67635
rect 74861 67589 74907 67635
rect 74985 67589 75031 67635
rect 75109 67589 75155 67635
rect 75233 67589 75279 67635
rect 75357 67589 75403 67635
rect 75481 67589 75527 67635
rect 75605 67589 75651 67635
rect 75729 67589 75775 67635
rect 75853 67589 75899 67635
rect 75977 67589 76023 67635
rect 76101 67589 76147 67635
rect 76225 67589 76271 67635
rect 76349 67589 76395 67635
rect 76473 67589 76519 67635
rect 76597 67589 76643 67635
rect 76721 67589 76767 67635
rect 76845 67589 76891 67635
rect 76969 67589 77015 67635
rect 77093 67589 77139 67635
rect 77217 67589 77263 67635
rect 77341 67589 77387 67635
rect 77465 67589 77511 67635
rect 77589 67589 77635 67635
rect 77713 67589 77759 67635
rect 77837 67589 77883 67635
rect 77961 67589 78007 67635
rect 78085 67589 78131 67635
rect 78209 67589 78255 67635
rect 78333 67589 78379 67635
rect 78457 67589 78503 67635
rect 78581 67589 78627 67635
rect 78705 67589 78751 67635
rect 78829 67589 78875 67635
rect 78953 67589 78999 67635
rect 79077 67589 79123 67635
rect 79201 67589 79247 67635
rect 79325 67589 79371 67635
rect 79449 67589 79495 67635
rect 79573 67589 79619 67635
rect 79697 67589 79743 67635
rect 79821 67589 79867 67635
rect 79945 67589 79991 67635
rect 80069 67589 80115 67635
rect 80193 67589 80239 67635
rect 80317 67589 80363 67635
rect 80441 67589 80487 67635
rect 80565 67589 80611 67635
rect 80689 67589 80735 67635
rect 80813 67589 80859 67635
rect 80937 67589 80983 67635
rect 81061 67589 81107 67635
rect 81185 67589 81231 67635
rect 81309 67589 81355 67635
rect 81433 67589 81479 67635
rect 81557 67589 81603 67635
rect 81681 67589 81727 67635
rect 81805 67589 81851 67635
rect 81929 67589 81975 67635
rect 82053 67589 82099 67635
rect 82177 67589 82223 67635
rect 82301 67589 82347 67635
rect 82425 67589 82471 67635
rect 82549 67589 82595 67635
rect 82673 67589 82719 67635
rect 82797 67589 82843 67635
rect 82921 67589 82967 67635
rect 83045 67589 83091 67635
rect 83169 67589 83215 67635
rect 83293 67589 83339 67635
rect 83417 67589 83463 67635
rect 83541 67589 83587 67635
rect 83665 67589 83711 67635
rect 83789 67589 83835 67635
rect 83913 67589 83959 67635
rect 84037 67589 84083 67635
rect 84161 67589 84207 67635
rect 84285 67589 84331 67635
rect 84409 67589 84455 67635
rect 84533 67589 84579 67635
rect 84657 67589 84703 67635
rect 84781 67589 84827 67635
rect 84905 67589 84951 67635
rect 85029 67589 85075 67635
rect 85153 67589 85199 67635
rect 85277 67589 85323 67635
rect 85401 67589 85447 67635
rect 85525 67589 85571 67635
rect 85649 67589 85695 67635
rect 89 67465 135 67511
rect 213 67465 259 67511
rect 337 67465 383 67511
rect 461 67465 507 67511
rect 585 67465 631 67511
rect 709 67465 755 67511
rect 833 67465 879 67511
rect 957 67465 1003 67511
rect 1081 67465 1127 67511
rect 1205 67465 1251 67511
rect 1329 67465 1375 67511
rect 1453 67465 1499 67511
rect 1577 67465 1623 67511
rect 1701 67465 1747 67511
rect 1825 67465 1871 67511
rect 1949 67465 1995 67511
rect 2073 67465 2119 67511
rect 2197 67465 2243 67511
rect 2321 67465 2367 67511
rect 2445 67465 2491 67511
rect 2569 67465 2615 67511
rect 2693 67465 2739 67511
rect 2817 67465 2863 67511
rect 2941 67465 2987 67511
rect 3065 67465 3111 67511
rect 3189 67465 3235 67511
rect 3313 67465 3359 67511
rect 3437 67465 3483 67511
rect 3561 67465 3607 67511
rect 3685 67465 3731 67511
rect 3809 67465 3855 67511
rect 3933 67465 3979 67511
rect 4057 67465 4103 67511
rect 4181 67465 4227 67511
rect 4305 67465 4351 67511
rect 4429 67465 4475 67511
rect 4553 67465 4599 67511
rect 4677 67465 4723 67511
rect 4801 67465 4847 67511
rect 4925 67465 4971 67511
rect 5049 67465 5095 67511
rect 5173 67465 5219 67511
rect 5297 67465 5343 67511
rect 5421 67465 5467 67511
rect 5545 67465 5591 67511
rect 5669 67465 5715 67511
rect 5793 67465 5839 67511
rect 5917 67465 5963 67511
rect 6041 67465 6087 67511
rect 6165 67465 6211 67511
rect 6289 67465 6335 67511
rect 6413 67465 6459 67511
rect 6537 67465 6583 67511
rect 6661 67465 6707 67511
rect 6785 67465 6831 67511
rect 6909 67465 6955 67511
rect 7033 67465 7079 67511
rect 7157 67465 7203 67511
rect 7281 67465 7327 67511
rect 7405 67465 7451 67511
rect 7529 67465 7575 67511
rect 7653 67465 7699 67511
rect 7777 67465 7823 67511
rect 7901 67465 7947 67511
rect 8025 67465 8071 67511
rect 8149 67465 8195 67511
rect 8273 67465 8319 67511
rect 8397 67465 8443 67511
rect 8521 67465 8567 67511
rect 8645 67465 8691 67511
rect 8769 67465 8815 67511
rect 8893 67465 8939 67511
rect 9017 67465 9063 67511
rect 9141 67465 9187 67511
rect 9265 67465 9311 67511
rect 9389 67465 9435 67511
rect 9513 67465 9559 67511
rect 9637 67465 9683 67511
rect 9761 67465 9807 67511
rect 9885 67465 9931 67511
rect 10009 67465 10055 67511
rect 10133 67465 10179 67511
rect 10257 67465 10303 67511
rect 10381 67465 10427 67511
rect 10505 67465 10551 67511
rect 10629 67465 10675 67511
rect 10753 67465 10799 67511
rect 10877 67465 10923 67511
rect 11001 67465 11047 67511
rect 11125 67465 11171 67511
rect 11249 67465 11295 67511
rect 11373 67465 11419 67511
rect 11497 67465 11543 67511
rect 11621 67465 11667 67511
rect 11745 67465 11791 67511
rect 11869 67465 11915 67511
rect 11993 67465 12039 67511
rect 12117 67465 12163 67511
rect 12241 67465 12287 67511
rect 12365 67465 12411 67511
rect 12489 67465 12535 67511
rect 12613 67465 12659 67511
rect 12737 67465 12783 67511
rect 12861 67465 12907 67511
rect 12985 67465 13031 67511
rect 13109 67465 13155 67511
rect 13233 67465 13279 67511
rect 13357 67465 13403 67511
rect 13481 67465 13527 67511
rect 13605 67465 13651 67511
rect 13729 67465 13775 67511
rect 13853 67465 13899 67511
rect 13977 67465 14023 67511
rect 14101 67465 14147 67511
rect 14225 67465 14271 67511
rect 14349 67465 14395 67511
rect 14473 67465 14519 67511
rect 14597 67465 14643 67511
rect 14721 67465 14767 67511
rect 14845 67465 14891 67511
rect 14969 67465 15015 67511
rect 15093 67465 15139 67511
rect 15217 67465 15263 67511
rect 15341 67465 15387 67511
rect 15465 67465 15511 67511
rect 15589 67465 15635 67511
rect 15713 67465 15759 67511
rect 15837 67465 15883 67511
rect 15961 67465 16007 67511
rect 16085 67465 16131 67511
rect 16209 67465 16255 67511
rect 16333 67465 16379 67511
rect 16457 67465 16503 67511
rect 16581 67465 16627 67511
rect 16705 67465 16751 67511
rect 16829 67465 16875 67511
rect 16953 67465 16999 67511
rect 17077 67465 17123 67511
rect 17201 67465 17247 67511
rect 17325 67465 17371 67511
rect 17449 67465 17495 67511
rect 17573 67465 17619 67511
rect 17697 67465 17743 67511
rect 17821 67465 17867 67511
rect 17945 67465 17991 67511
rect 18069 67465 18115 67511
rect 18193 67465 18239 67511
rect 18317 67465 18363 67511
rect 18441 67465 18487 67511
rect 18565 67465 18611 67511
rect 18689 67465 18735 67511
rect 18813 67465 18859 67511
rect 18937 67465 18983 67511
rect 19061 67465 19107 67511
rect 19185 67465 19231 67511
rect 19309 67465 19355 67511
rect 19433 67465 19479 67511
rect 19557 67465 19603 67511
rect 19681 67465 19727 67511
rect 19805 67465 19851 67511
rect 19929 67465 19975 67511
rect 20053 67465 20099 67511
rect 20177 67465 20223 67511
rect 20301 67465 20347 67511
rect 20425 67465 20471 67511
rect 20549 67465 20595 67511
rect 20673 67465 20719 67511
rect 20797 67465 20843 67511
rect 20921 67465 20967 67511
rect 21045 67465 21091 67511
rect 21169 67465 21215 67511
rect 21293 67465 21339 67511
rect 21417 67465 21463 67511
rect 21541 67465 21587 67511
rect 21665 67465 21711 67511
rect 21789 67465 21835 67511
rect 21913 67465 21959 67511
rect 22037 67465 22083 67511
rect 22161 67465 22207 67511
rect 22285 67465 22331 67511
rect 22409 67465 22455 67511
rect 22533 67465 22579 67511
rect 22657 67465 22703 67511
rect 22781 67465 22827 67511
rect 22905 67465 22951 67511
rect 23029 67465 23075 67511
rect 23153 67465 23199 67511
rect 23277 67465 23323 67511
rect 23401 67465 23447 67511
rect 23525 67465 23571 67511
rect 23649 67465 23695 67511
rect 23773 67465 23819 67511
rect 23897 67465 23943 67511
rect 24021 67465 24067 67511
rect 24145 67465 24191 67511
rect 24269 67465 24315 67511
rect 24393 67465 24439 67511
rect 24517 67465 24563 67511
rect 24641 67465 24687 67511
rect 24765 67465 24811 67511
rect 24889 67465 24935 67511
rect 25013 67465 25059 67511
rect 25137 67465 25183 67511
rect 25261 67465 25307 67511
rect 25385 67465 25431 67511
rect 25509 67465 25555 67511
rect 25633 67465 25679 67511
rect 25757 67465 25803 67511
rect 25881 67465 25927 67511
rect 26005 67465 26051 67511
rect 26129 67465 26175 67511
rect 26253 67465 26299 67511
rect 26377 67465 26423 67511
rect 26501 67465 26547 67511
rect 26625 67465 26671 67511
rect 26749 67465 26795 67511
rect 26873 67465 26919 67511
rect 26997 67465 27043 67511
rect 27121 67465 27167 67511
rect 27245 67465 27291 67511
rect 27369 67465 27415 67511
rect 27493 67465 27539 67511
rect 27617 67465 27663 67511
rect 27741 67465 27787 67511
rect 27865 67465 27911 67511
rect 27989 67465 28035 67511
rect 28113 67465 28159 67511
rect 28237 67465 28283 67511
rect 28361 67465 28407 67511
rect 28485 67465 28531 67511
rect 28609 67465 28655 67511
rect 28733 67465 28779 67511
rect 28857 67465 28903 67511
rect 28981 67465 29027 67511
rect 29105 67465 29151 67511
rect 29229 67465 29275 67511
rect 29353 67465 29399 67511
rect 29477 67465 29523 67511
rect 29601 67465 29647 67511
rect 29725 67465 29771 67511
rect 29849 67465 29895 67511
rect 29973 67465 30019 67511
rect 30097 67465 30143 67511
rect 30221 67465 30267 67511
rect 30345 67465 30391 67511
rect 30469 67465 30515 67511
rect 30593 67465 30639 67511
rect 30717 67465 30763 67511
rect 30841 67465 30887 67511
rect 30965 67465 31011 67511
rect 31089 67465 31135 67511
rect 31213 67465 31259 67511
rect 31337 67465 31383 67511
rect 31461 67465 31507 67511
rect 31585 67465 31631 67511
rect 31709 67465 31755 67511
rect 31833 67465 31879 67511
rect 31957 67465 32003 67511
rect 32081 67465 32127 67511
rect 32205 67465 32251 67511
rect 32329 67465 32375 67511
rect 32453 67465 32499 67511
rect 32577 67465 32623 67511
rect 32701 67465 32747 67511
rect 32825 67465 32871 67511
rect 32949 67465 32995 67511
rect 33073 67465 33119 67511
rect 33197 67465 33243 67511
rect 33321 67465 33367 67511
rect 33445 67465 33491 67511
rect 33569 67465 33615 67511
rect 33693 67465 33739 67511
rect 33817 67465 33863 67511
rect 33941 67465 33987 67511
rect 34065 67465 34111 67511
rect 34189 67465 34235 67511
rect 34313 67465 34359 67511
rect 34437 67465 34483 67511
rect 34561 67465 34607 67511
rect 34685 67465 34731 67511
rect 34809 67465 34855 67511
rect 34933 67465 34979 67511
rect 35057 67465 35103 67511
rect 35181 67465 35227 67511
rect 35305 67465 35351 67511
rect 35429 67465 35475 67511
rect 35553 67465 35599 67511
rect 35677 67465 35723 67511
rect 35801 67465 35847 67511
rect 35925 67465 35971 67511
rect 36049 67465 36095 67511
rect 36173 67465 36219 67511
rect 36297 67465 36343 67511
rect 36421 67465 36467 67511
rect 36545 67465 36591 67511
rect 36669 67465 36715 67511
rect 36793 67465 36839 67511
rect 36917 67465 36963 67511
rect 37041 67465 37087 67511
rect 37165 67465 37211 67511
rect 37289 67465 37335 67511
rect 37413 67465 37459 67511
rect 37537 67465 37583 67511
rect 37661 67465 37707 67511
rect 37785 67465 37831 67511
rect 37909 67465 37955 67511
rect 38033 67465 38079 67511
rect 38157 67465 38203 67511
rect 38281 67465 38327 67511
rect 38405 67465 38451 67511
rect 38529 67465 38575 67511
rect 38653 67465 38699 67511
rect 38777 67465 38823 67511
rect 38901 67465 38947 67511
rect 39025 67465 39071 67511
rect 39149 67465 39195 67511
rect 39273 67465 39319 67511
rect 39397 67465 39443 67511
rect 39521 67465 39567 67511
rect 39645 67465 39691 67511
rect 39769 67465 39815 67511
rect 39893 67465 39939 67511
rect 40017 67465 40063 67511
rect 40141 67465 40187 67511
rect 40265 67465 40311 67511
rect 40389 67465 40435 67511
rect 40513 67465 40559 67511
rect 40637 67465 40683 67511
rect 40761 67465 40807 67511
rect 40885 67465 40931 67511
rect 41009 67465 41055 67511
rect 41133 67465 41179 67511
rect 41257 67465 41303 67511
rect 41381 67465 41427 67511
rect 41505 67465 41551 67511
rect 41629 67465 41675 67511
rect 41753 67465 41799 67511
rect 41877 67465 41923 67511
rect 42001 67465 42047 67511
rect 42125 67465 42171 67511
rect 42249 67465 42295 67511
rect 42373 67465 42419 67511
rect 42497 67465 42543 67511
rect 42621 67465 42667 67511
rect 42745 67465 42791 67511
rect 42869 67465 42915 67511
rect 42993 67465 43039 67511
rect 43117 67465 43163 67511
rect 43241 67465 43287 67511
rect 43365 67465 43411 67511
rect 43489 67465 43535 67511
rect 43613 67465 43659 67511
rect 43737 67465 43783 67511
rect 43861 67465 43907 67511
rect 43985 67465 44031 67511
rect 44109 67465 44155 67511
rect 44233 67465 44279 67511
rect 44357 67465 44403 67511
rect 44481 67465 44527 67511
rect 44605 67465 44651 67511
rect 44729 67465 44775 67511
rect 44853 67465 44899 67511
rect 44977 67465 45023 67511
rect 45101 67465 45147 67511
rect 45225 67465 45271 67511
rect 45349 67465 45395 67511
rect 45473 67465 45519 67511
rect 45597 67465 45643 67511
rect 45721 67465 45767 67511
rect 45845 67465 45891 67511
rect 45969 67465 46015 67511
rect 46093 67465 46139 67511
rect 46217 67465 46263 67511
rect 46341 67465 46387 67511
rect 46465 67465 46511 67511
rect 46589 67465 46635 67511
rect 46713 67465 46759 67511
rect 46837 67465 46883 67511
rect 46961 67465 47007 67511
rect 47085 67465 47131 67511
rect 47209 67465 47255 67511
rect 47333 67465 47379 67511
rect 47457 67465 47503 67511
rect 47581 67465 47627 67511
rect 47705 67465 47751 67511
rect 47829 67465 47875 67511
rect 47953 67465 47999 67511
rect 48077 67465 48123 67511
rect 48201 67465 48247 67511
rect 48325 67465 48371 67511
rect 48449 67465 48495 67511
rect 48573 67465 48619 67511
rect 48697 67465 48743 67511
rect 48821 67465 48867 67511
rect 48945 67465 48991 67511
rect 49069 67465 49115 67511
rect 49193 67465 49239 67511
rect 49317 67465 49363 67511
rect 49441 67465 49487 67511
rect 49565 67465 49611 67511
rect 49689 67465 49735 67511
rect 49813 67465 49859 67511
rect 49937 67465 49983 67511
rect 50061 67465 50107 67511
rect 50185 67465 50231 67511
rect 50309 67465 50355 67511
rect 50433 67465 50479 67511
rect 50557 67465 50603 67511
rect 50681 67465 50727 67511
rect 50805 67465 50851 67511
rect 50929 67465 50975 67511
rect 51053 67465 51099 67511
rect 51177 67465 51223 67511
rect 51301 67465 51347 67511
rect 51425 67465 51471 67511
rect 51549 67465 51595 67511
rect 51673 67465 51719 67511
rect 51797 67465 51843 67511
rect 51921 67465 51967 67511
rect 52045 67465 52091 67511
rect 52169 67465 52215 67511
rect 52293 67465 52339 67511
rect 52417 67465 52463 67511
rect 52541 67465 52587 67511
rect 52665 67465 52711 67511
rect 52789 67465 52835 67511
rect 52913 67465 52959 67511
rect 53037 67465 53083 67511
rect 53161 67465 53207 67511
rect 53285 67465 53331 67511
rect 53409 67465 53455 67511
rect 53533 67465 53579 67511
rect 53657 67465 53703 67511
rect 53781 67465 53827 67511
rect 53905 67465 53951 67511
rect 54029 67465 54075 67511
rect 54153 67465 54199 67511
rect 54277 67465 54323 67511
rect 54401 67465 54447 67511
rect 54525 67465 54571 67511
rect 54649 67465 54695 67511
rect 54773 67465 54819 67511
rect 54897 67465 54943 67511
rect 55021 67465 55067 67511
rect 55145 67465 55191 67511
rect 55269 67465 55315 67511
rect 55393 67465 55439 67511
rect 55517 67465 55563 67511
rect 55641 67465 55687 67511
rect 55765 67465 55811 67511
rect 55889 67465 55935 67511
rect 56013 67465 56059 67511
rect 56137 67465 56183 67511
rect 56261 67465 56307 67511
rect 56385 67465 56431 67511
rect 56509 67465 56555 67511
rect 56633 67465 56679 67511
rect 56757 67465 56803 67511
rect 56881 67465 56927 67511
rect 57005 67465 57051 67511
rect 57129 67465 57175 67511
rect 57253 67465 57299 67511
rect 57377 67465 57423 67511
rect 57501 67465 57547 67511
rect 57625 67465 57671 67511
rect 57749 67465 57795 67511
rect 57873 67465 57919 67511
rect 57997 67465 58043 67511
rect 58121 67465 58167 67511
rect 58245 67465 58291 67511
rect 58369 67465 58415 67511
rect 58493 67465 58539 67511
rect 58617 67465 58663 67511
rect 58741 67465 58787 67511
rect 58865 67465 58911 67511
rect 58989 67465 59035 67511
rect 59113 67465 59159 67511
rect 59237 67465 59283 67511
rect 59361 67465 59407 67511
rect 59485 67465 59531 67511
rect 59609 67465 59655 67511
rect 59733 67465 59779 67511
rect 59857 67465 59903 67511
rect 59981 67465 60027 67511
rect 60105 67465 60151 67511
rect 60229 67465 60275 67511
rect 60353 67465 60399 67511
rect 60477 67465 60523 67511
rect 60601 67465 60647 67511
rect 60725 67465 60771 67511
rect 60849 67465 60895 67511
rect 60973 67465 61019 67511
rect 61097 67465 61143 67511
rect 61221 67465 61267 67511
rect 61345 67465 61391 67511
rect 61469 67465 61515 67511
rect 61593 67465 61639 67511
rect 61717 67465 61763 67511
rect 61841 67465 61887 67511
rect 61965 67465 62011 67511
rect 62089 67465 62135 67511
rect 62213 67465 62259 67511
rect 62337 67465 62383 67511
rect 62461 67465 62507 67511
rect 62585 67465 62631 67511
rect 62709 67465 62755 67511
rect 62833 67465 62879 67511
rect 62957 67465 63003 67511
rect 63081 67465 63127 67511
rect 63205 67465 63251 67511
rect 63329 67465 63375 67511
rect 63453 67465 63499 67511
rect 63577 67465 63623 67511
rect 63701 67465 63747 67511
rect 63825 67465 63871 67511
rect 63949 67465 63995 67511
rect 64073 67465 64119 67511
rect 64197 67465 64243 67511
rect 64321 67465 64367 67511
rect 64445 67465 64491 67511
rect 64569 67465 64615 67511
rect 64693 67465 64739 67511
rect 64817 67465 64863 67511
rect 64941 67465 64987 67511
rect 65065 67465 65111 67511
rect 65189 67465 65235 67511
rect 65313 67465 65359 67511
rect 65437 67465 65483 67511
rect 65561 67465 65607 67511
rect 65685 67465 65731 67511
rect 65809 67465 65855 67511
rect 65933 67465 65979 67511
rect 66057 67465 66103 67511
rect 66181 67465 66227 67511
rect 66305 67465 66351 67511
rect 66429 67465 66475 67511
rect 66553 67465 66599 67511
rect 66677 67465 66723 67511
rect 66801 67465 66847 67511
rect 66925 67465 66971 67511
rect 67049 67465 67095 67511
rect 67173 67465 67219 67511
rect 67297 67465 67343 67511
rect 67421 67465 67467 67511
rect 67545 67465 67591 67511
rect 67669 67465 67715 67511
rect 67793 67465 67839 67511
rect 67917 67465 67963 67511
rect 68041 67465 68087 67511
rect 68165 67465 68211 67511
rect 68289 67465 68335 67511
rect 68413 67465 68459 67511
rect 68537 67465 68583 67511
rect 68661 67465 68707 67511
rect 68785 67465 68831 67511
rect 68909 67465 68955 67511
rect 69033 67465 69079 67511
rect 69157 67465 69203 67511
rect 69281 67465 69327 67511
rect 69405 67465 69451 67511
rect 69529 67465 69575 67511
rect 69653 67465 69699 67511
rect 69777 67465 69823 67511
rect 69901 67465 69947 67511
rect 70025 67465 70071 67511
rect 70149 67465 70195 67511
rect 70273 67465 70319 67511
rect 70397 67465 70443 67511
rect 70521 67465 70567 67511
rect 70645 67465 70691 67511
rect 70769 67465 70815 67511
rect 70893 67465 70939 67511
rect 71017 67465 71063 67511
rect 71141 67465 71187 67511
rect 71265 67465 71311 67511
rect 71389 67465 71435 67511
rect 71513 67465 71559 67511
rect 71637 67465 71683 67511
rect 71761 67465 71807 67511
rect 71885 67465 71931 67511
rect 72009 67465 72055 67511
rect 72133 67465 72179 67511
rect 72257 67465 72303 67511
rect 72381 67465 72427 67511
rect 72505 67465 72551 67511
rect 72629 67465 72675 67511
rect 72753 67465 72799 67511
rect 72877 67465 72923 67511
rect 73001 67465 73047 67511
rect 73125 67465 73171 67511
rect 73249 67465 73295 67511
rect 73373 67465 73419 67511
rect 73497 67465 73543 67511
rect 73621 67465 73667 67511
rect 73745 67465 73791 67511
rect 73869 67465 73915 67511
rect 73993 67465 74039 67511
rect 74117 67465 74163 67511
rect 74241 67465 74287 67511
rect 74365 67465 74411 67511
rect 74489 67465 74535 67511
rect 74613 67465 74659 67511
rect 74737 67465 74783 67511
rect 74861 67465 74907 67511
rect 74985 67465 75031 67511
rect 75109 67465 75155 67511
rect 75233 67465 75279 67511
rect 75357 67465 75403 67511
rect 75481 67465 75527 67511
rect 75605 67465 75651 67511
rect 75729 67465 75775 67511
rect 75853 67465 75899 67511
rect 75977 67465 76023 67511
rect 76101 67465 76147 67511
rect 76225 67465 76271 67511
rect 76349 67465 76395 67511
rect 76473 67465 76519 67511
rect 76597 67465 76643 67511
rect 76721 67465 76767 67511
rect 76845 67465 76891 67511
rect 76969 67465 77015 67511
rect 77093 67465 77139 67511
rect 77217 67465 77263 67511
rect 77341 67465 77387 67511
rect 77465 67465 77511 67511
rect 77589 67465 77635 67511
rect 77713 67465 77759 67511
rect 77837 67465 77883 67511
rect 77961 67465 78007 67511
rect 78085 67465 78131 67511
rect 78209 67465 78255 67511
rect 78333 67465 78379 67511
rect 78457 67465 78503 67511
rect 78581 67465 78627 67511
rect 78705 67465 78751 67511
rect 78829 67465 78875 67511
rect 78953 67465 78999 67511
rect 79077 67465 79123 67511
rect 79201 67465 79247 67511
rect 79325 67465 79371 67511
rect 79449 67465 79495 67511
rect 79573 67465 79619 67511
rect 79697 67465 79743 67511
rect 79821 67465 79867 67511
rect 79945 67465 79991 67511
rect 80069 67465 80115 67511
rect 80193 67465 80239 67511
rect 80317 67465 80363 67511
rect 80441 67465 80487 67511
rect 80565 67465 80611 67511
rect 80689 67465 80735 67511
rect 80813 67465 80859 67511
rect 80937 67465 80983 67511
rect 81061 67465 81107 67511
rect 81185 67465 81231 67511
rect 81309 67465 81355 67511
rect 81433 67465 81479 67511
rect 81557 67465 81603 67511
rect 81681 67465 81727 67511
rect 81805 67465 81851 67511
rect 81929 67465 81975 67511
rect 82053 67465 82099 67511
rect 82177 67465 82223 67511
rect 82301 67465 82347 67511
rect 82425 67465 82471 67511
rect 82549 67465 82595 67511
rect 82673 67465 82719 67511
rect 82797 67465 82843 67511
rect 82921 67465 82967 67511
rect 83045 67465 83091 67511
rect 83169 67465 83215 67511
rect 83293 67465 83339 67511
rect 83417 67465 83463 67511
rect 83541 67465 83587 67511
rect 83665 67465 83711 67511
rect 83789 67465 83835 67511
rect 83913 67465 83959 67511
rect 84037 67465 84083 67511
rect 84161 67465 84207 67511
rect 84285 67465 84331 67511
rect 84409 67465 84455 67511
rect 84533 67465 84579 67511
rect 84657 67465 84703 67511
rect 84781 67465 84827 67511
rect 84905 67465 84951 67511
rect 85029 67465 85075 67511
rect 85153 67465 85199 67511
rect 85277 67465 85323 67511
rect 85401 67465 85447 67511
rect 85525 67465 85571 67511
rect 85649 67465 85695 67511
rect 89 1117 435 67363
rect 27116 1117 27462 67363
rect 27564 35996 28410 67342
rect 56110 35996 56956 67342
rect 27564 34242 56910 34588
rect 57024 1117 57370 67363
rect 85451 1117 85797 67363
rect 89 969 135 1015
rect 213 969 259 1015
rect 337 969 383 1015
rect 461 969 507 1015
rect 585 969 631 1015
rect 709 969 755 1015
rect 833 969 879 1015
rect 957 969 1003 1015
rect 1081 969 1127 1015
rect 1205 969 1251 1015
rect 1329 969 1375 1015
rect 1453 969 1499 1015
rect 1577 969 1623 1015
rect 1701 969 1747 1015
rect 1825 969 1871 1015
rect 1949 969 1995 1015
rect 2073 969 2119 1015
rect 2197 969 2243 1015
rect 2321 969 2367 1015
rect 2445 969 2491 1015
rect 2569 969 2615 1015
rect 2693 969 2739 1015
rect 2817 969 2863 1015
rect 2941 969 2987 1015
rect 3065 969 3111 1015
rect 3189 969 3235 1015
rect 3313 969 3359 1015
rect 3437 969 3483 1015
rect 3561 969 3607 1015
rect 3685 969 3731 1015
rect 3809 969 3855 1015
rect 3933 969 3979 1015
rect 4057 969 4103 1015
rect 4181 969 4227 1015
rect 4305 969 4351 1015
rect 4429 969 4475 1015
rect 4553 969 4599 1015
rect 4677 969 4723 1015
rect 4801 969 4847 1015
rect 4925 969 4971 1015
rect 5049 969 5095 1015
rect 5173 969 5219 1015
rect 5297 969 5343 1015
rect 5421 969 5467 1015
rect 5545 969 5591 1015
rect 5669 969 5715 1015
rect 5793 969 5839 1015
rect 5917 969 5963 1015
rect 6041 969 6087 1015
rect 6165 969 6211 1015
rect 6289 969 6335 1015
rect 6413 969 6459 1015
rect 6537 969 6583 1015
rect 6661 969 6707 1015
rect 6785 969 6831 1015
rect 6909 969 6955 1015
rect 7033 969 7079 1015
rect 7157 969 7203 1015
rect 7281 969 7327 1015
rect 7405 969 7451 1015
rect 7529 969 7575 1015
rect 7653 969 7699 1015
rect 7777 969 7823 1015
rect 7901 969 7947 1015
rect 8025 969 8071 1015
rect 8149 969 8195 1015
rect 8273 969 8319 1015
rect 8397 969 8443 1015
rect 8521 969 8567 1015
rect 8645 969 8691 1015
rect 8769 969 8815 1015
rect 8893 969 8939 1015
rect 9017 969 9063 1015
rect 9141 969 9187 1015
rect 9265 969 9311 1015
rect 9389 969 9435 1015
rect 9513 969 9559 1015
rect 9637 969 9683 1015
rect 9761 969 9807 1015
rect 9885 969 9931 1015
rect 10009 969 10055 1015
rect 10133 969 10179 1015
rect 10257 969 10303 1015
rect 10381 969 10427 1015
rect 10505 969 10551 1015
rect 10629 969 10675 1015
rect 10753 969 10799 1015
rect 10877 969 10923 1015
rect 11001 969 11047 1015
rect 11125 969 11171 1015
rect 11249 969 11295 1015
rect 11373 969 11419 1015
rect 11497 969 11543 1015
rect 11621 969 11667 1015
rect 11745 969 11791 1015
rect 11869 969 11915 1015
rect 11993 969 12039 1015
rect 12117 969 12163 1015
rect 12241 969 12287 1015
rect 12365 969 12411 1015
rect 12489 969 12535 1015
rect 12613 969 12659 1015
rect 12737 969 12783 1015
rect 12861 969 12907 1015
rect 12985 969 13031 1015
rect 13109 969 13155 1015
rect 13233 969 13279 1015
rect 13357 969 13403 1015
rect 13481 969 13527 1015
rect 13605 969 13651 1015
rect 13729 969 13775 1015
rect 13853 969 13899 1015
rect 13977 969 14023 1015
rect 14101 969 14147 1015
rect 14225 969 14271 1015
rect 14349 969 14395 1015
rect 14473 969 14519 1015
rect 14597 969 14643 1015
rect 14721 969 14767 1015
rect 14845 969 14891 1015
rect 14969 969 15015 1015
rect 15093 969 15139 1015
rect 15217 969 15263 1015
rect 15341 969 15387 1015
rect 15465 969 15511 1015
rect 15589 969 15635 1015
rect 15713 969 15759 1015
rect 15837 969 15883 1015
rect 15961 969 16007 1015
rect 16085 969 16131 1015
rect 16209 969 16255 1015
rect 16333 969 16379 1015
rect 16457 969 16503 1015
rect 16581 969 16627 1015
rect 16705 969 16751 1015
rect 16829 969 16875 1015
rect 16953 969 16999 1015
rect 17077 969 17123 1015
rect 17201 969 17247 1015
rect 17325 969 17371 1015
rect 17449 969 17495 1015
rect 17573 969 17619 1015
rect 17697 969 17743 1015
rect 17821 969 17867 1015
rect 17945 969 17991 1015
rect 18069 969 18115 1015
rect 18193 969 18239 1015
rect 18317 969 18363 1015
rect 18441 969 18487 1015
rect 18565 969 18611 1015
rect 18689 969 18735 1015
rect 18813 969 18859 1015
rect 18937 969 18983 1015
rect 19061 969 19107 1015
rect 19185 969 19231 1015
rect 19309 969 19355 1015
rect 19433 969 19479 1015
rect 19557 969 19603 1015
rect 19681 969 19727 1015
rect 19805 969 19851 1015
rect 19929 969 19975 1015
rect 20053 969 20099 1015
rect 20177 969 20223 1015
rect 20301 969 20347 1015
rect 20425 969 20471 1015
rect 20549 969 20595 1015
rect 20673 969 20719 1015
rect 20797 969 20843 1015
rect 20921 969 20967 1015
rect 21045 969 21091 1015
rect 21169 969 21215 1015
rect 21293 969 21339 1015
rect 21417 969 21463 1015
rect 21541 969 21587 1015
rect 21665 969 21711 1015
rect 21789 969 21835 1015
rect 21913 969 21959 1015
rect 22037 969 22083 1015
rect 22161 969 22207 1015
rect 22285 969 22331 1015
rect 22409 969 22455 1015
rect 22533 969 22579 1015
rect 22657 969 22703 1015
rect 22781 969 22827 1015
rect 22905 969 22951 1015
rect 23029 969 23075 1015
rect 23153 969 23199 1015
rect 23277 969 23323 1015
rect 23401 969 23447 1015
rect 23525 969 23571 1015
rect 23649 969 23695 1015
rect 23773 969 23819 1015
rect 23897 969 23943 1015
rect 24021 969 24067 1015
rect 24145 969 24191 1015
rect 24269 969 24315 1015
rect 24393 969 24439 1015
rect 24517 969 24563 1015
rect 24641 969 24687 1015
rect 24765 969 24811 1015
rect 24889 969 24935 1015
rect 25013 969 25059 1015
rect 25137 969 25183 1015
rect 25261 969 25307 1015
rect 25385 969 25431 1015
rect 25509 969 25555 1015
rect 25633 969 25679 1015
rect 25757 969 25803 1015
rect 25881 969 25927 1015
rect 26005 969 26051 1015
rect 26129 969 26175 1015
rect 26253 969 26299 1015
rect 26377 969 26423 1015
rect 26501 969 26547 1015
rect 26625 969 26671 1015
rect 26749 969 26795 1015
rect 26873 969 26919 1015
rect 26997 969 27043 1015
rect 27121 969 27167 1015
rect 27245 969 27291 1015
rect 27369 969 27415 1015
rect 27493 969 27539 1015
rect 27617 969 27663 1015
rect 27741 969 27787 1015
rect 27865 969 27911 1015
rect 27989 969 28035 1015
rect 28113 969 28159 1015
rect 28237 969 28283 1015
rect 28361 969 28407 1015
rect 28485 969 28531 1015
rect 28609 969 28655 1015
rect 28733 969 28779 1015
rect 28857 969 28903 1015
rect 28981 969 29027 1015
rect 29105 969 29151 1015
rect 29229 969 29275 1015
rect 29353 969 29399 1015
rect 29477 969 29523 1015
rect 29601 969 29647 1015
rect 29725 969 29771 1015
rect 29849 969 29895 1015
rect 29973 969 30019 1015
rect 30097 969 30143 1015
rect 30221 969 30267 1015
rect 30345 969 30391 1015
rect 30469 969 30515 1015
rect 30593 969 30639 1015
rect 30717 969 30763 1015
rect 30841 969 30887 1015
rect 30965 969 31011 1015
rect 31089 969 31135 1015
rect 31213 969 31259 1015
rect 31337 969 31383 1015
rect 31461 969 31507 1015
rect 31585 969 31631 1015
rect 31709 969 31755 1015
rect 31833 969 31879 1015
rect 31957 969 32003 1015
rect 32081 969 32127 1015
rect 32205 969 32251 1015
rect 32329 969 32375 1015
rect 32453 969 32499 1015
rect 32577 969 32623 1015
rect 32701 969 32747 1015
rect 32825 969 32871 1015
rect 32949 969 32995 1015
rect 33073 969 33119 1015
rect 33197 969 33243 1015
rect 33321 969 33367 1015
rect 33445 969 33491 1015
rect 33569 969 33615 1015
rect 33693 969 33739 1015
rect 33817 969 33863 1015
rect 33941 969 33987 1015
rect 34065 969 34111 1015
rect 34189 969 34235 1015
rect 34313 969 34359 1015
rect 34437 969 34483 1015
rect 34561 969 34607 1015
rect 34685 969 34731 1015
rect 34809 969 34855 1015
rect 34933 969 34979 1015
rect 35057 969 35103 1015
rect 35181 969 35227 1015
rect 35305 969 35351 1015
rect 35429 969 35475 1015
rect 35553 969 35599 1015
rect 35677 969 35723 1015
rect 35801 969 35847 1015
rect 35925 969 35971 1015
rect 36049 969 36095 1015
rect 36173 969 36219 1015
rect 36297 969 36343 1015
rect 36421 969 36467 1015
rect 36545 969 36591 1015
rect 36669 969 36715 1015
rect 36793 969 36839 1015
rect 36917 969 36963 1015
rect 37041 969 37087 1015
rect 37165 969 37211 1015
rect 37289 969 37335 1015
rect 37413 969 37459 1015
rect 37537 969 37583 1015
rect 37661 969 37707 1015
rect 37785 969 37831 1015
rect 37909 969 37955 1015
rect 38033 969 38079 1015
rect 38157 969 38203 1015
rect 38281 969 38327 1015
rect 38405 969 38451 1015
rect 38529 969 38575 1015
rect 38653 969 38699 1015
rect 38777 969 38823 1015
rect 38901 969 38947 1015
rect 39025 969 39071 1015
rect 39149 969 39195 1015
rect 39273 969 39319 1015
rect 39397 969 39443 1015
rect 39521 969 39567 1015
rect 39645 969 39691 1015
rect 39769 969 39815 1015
rect 39893 969 39939 1015
rect 40017 969 40063 1015
rect 40141 969 40187 1015
rect 40265 969 40311 1015
rect 40389 969 40435 1015
rect 40513 969 40559 1015
rect 40637 969 40683 1015
rect 40761 969 40807 1015
rect 40885 969 40931 1015
rect 41009 969 41055 1015
rect 41133 969 41179 1015
rect 41257 969 41303 1015
rect 41381 969 41427 1015
rect 41505 969 41551 1015
rect 41629 969 41675 1015
rect 41753 969 41799 1015
rect 41877 969 41923 1015
rect 42001 969 42047 1015
rect 42125 969 42171 1015
rect 42249 969 42295 1015
rect 42373 969 42419 1015
rect 42497 969 42543 1015
rect 42621 969 42667 1015
rect 42745 969 42791 1015
rect 42869 969 42915 1015
rect 42993 969 43039 1015
rect 43117 969 43163 1015
rect 43241 969 43287 1015
rect 43365 969 43411 1015
rect 43489 969 43535 1015
rect 43613 969 43659 1015
rect 43737 969 43783 1015
rect 43861 969 43907 1015
rect 43985 969 44031 1015
rect 44109 969 44155 1015
rect 44233 969 44279 1015
rect 44357 969 44403 1015
rect 44481 969 44527 1015
rect 44605 969 44651 1015
rect 44729 969 44775 1015
rect 44853 969 44899 1015
rect 44977 969 45023 1015
rect 45101 969 45147 1015
rect 45225 969 45271 1015
rect 45349 969 45395 1015
rect 45473 969 45519 1015
rect 45597 969 45643 1015
rect 45721 969 45767 1015
rect 45845 969 45891 1015
rect 45969 969 46015 1015
rect 46093 969 46139 1015
rect 46217 969 46263 1015
rect 46341 969 46387 1015
rect 46465 969 46511 1015
rect 46589 969 46635 1015
rect 46713 969 46759 1015
rect 46837 969 46883 1015
rect 46961 969 47007 1015
rect 47085 969 47131 1015
rect 47209 969 47255 1015
rect 47333 969 47379 1015
rect 47457 969 47503 1015
rect 47581 969 47627 1015
rect 47705 969 47751 1015
rect 47829 969 47875 1015
rect 47953 969 47999 1015
rect 48077 969 48123 1015
rect 48201 969 48247 1015
rect 48325 969 48371 1015
rect 48449 969 48495 1015
rect 48573 969 48619 1015
rect 48697 969 48743 1015
rect 48821 969 48867 1015
rect 48945 969 48991 1015
rect 49069 969 49115 1015
rect 49193 969 49239 1015
rect 49317 969 49363 1015
rect 49441 969 49487 1015
rect 49565 969 49611 1015
rect 49689 969 49735 1015
rect 49813 969 49859 1015
rect 49937 969 49983 1015
rect 50061 969 50107 1015
rect 50185 969 50231 1015
rect 50309 969 50355 1015
rect 50433 969 50479 1015
rect 50557 969 50603 1015
rect 50681 969 50727 1015
rect 50805 969 50851 1015
rect 50929 969 50975 1015
rect 51053 969 51099 1015
rect 51177 969 51223 1015
rect 51301 969 51347 1015
rect 51425 969 51471 1015
rect 51549 969 51595 1015
rect 51673 969 51719 1015
rect 51797 969 51843 1015
rect 51921 969 51967 1015
rect 52045 969 52091 1015
rect 52169 969 52215 1015
rect 52293 969 52339 1015
rect 52417 969 52463 1015
rect 52541 969 52587 1015
rect 52665 969 52711 1015
rect 52789 969 52835 1015
rect 52913 969 52959 1015
rect 53037 969 53083 1015
rect 53161 969 53207 1015
rect 53285 969 53331 1015
rect 53409 969 53455 1015
rect 53533 969 53579 1015
rect 53657 969 53703 1015
rect 53781 969 53827 1015
rect 53905 969 53951 1015
rect 54029 969 54075 1015
rect 54153 969 54199 1015
rect 54277 969 54323 1015
rect 54401 969 54447 1015
rect 54525 969 54571 1015
rect 54649 969 54695 1015
rect 54773 969 54819 1015
rect 54897 969 54943 1015
rect 55021 969 55067 1015
rect 55145 969 55191 1015
rect 55269 969 55315 1015
rect 55393 969 55439 1015
rect 55517 969 55563 1015
rect 55641 969 55687 1015
rect 55765 969 55811 1015
rect 55889 969 55935 1015
rect 56013 969 56059 1015
rect 56137 969 56183 1015
rect 56261 969 56307 1015
rect 56385 969 56431 1015
rect 56509 969 56555 1015
rect 56633 969 56679 1015
rect 56757 969 56803 1015
rect 56881 969 56927 1015
rect 57005 969 57051 1015
rect 57129 969 57175 1015
rect 57253 969 57299 1015
rect 57377 969 57423 1015
rect 57501 969 57547 1015
rect 57625 969 57671 1015
rect 57749 969 57795 1015
rect 57873 969 57919 1015
rect 57997 969 58043 1015
rect 58121 969 58167 1015
rect 58245 969 58291 1015
rect 58369 969 58415 1015
rect 58493 969 58539 1015
rect 58617 969 58663 1015
rect 58741 969 58787 1015
rect 58865 969 58911 1015
rect 58989 969 59035 1015
rect 59113 969 59159 1015
rect 59237 969 59283 1015
rect 59361 969 59407 1015
rect 59485 969 59531 1015
rect 59609 969 59655 1015
rect 59733 969 59779 1015
rect 59857 969 59903 1015
rect 59981 969 60027 1015
rect 60105 969 60151 1015
rect 60229 969 60275 1015
rect 60353 969 60399 1015
rect 60477 969 60523 1015
rect 60601 969 60647 1015
rect 60725 969 60771 1015
rect 60849 969 60895 1015
rect 60973 969 61019 1015
rect 61097 969 61143 1015
rect 61221 969 61267 1015
rect 61345 969 61391 1015
rect 61469 969 61515 1015
rect 61593 969 61639 1015
rect 61717 969 61763 1015
rect 61841 969 61887 1015
rect 61965 969 62011 1015
rect 62089 969 62135 1015
rect 62213 969 62259 1015
rect 62337 969 62383 1015
rect 62461 969 62507 1015
rect 62585 969 62631 1015
rect 62709 969 62755 1015
rect 62833 969 62879 1015
rect 62957 969 63003 1015
rect 63081 969 63127 1015
rect 63205 969 63251 1015
rect 63329 969 63375 1015
rect 63453 969 63499 1015
rect 63577 969 63623 1015
rect 63701 969 63747 1015
rect 63825 969 63871 1015
rect 63949 969 63995 1015
rect 64073 969 64119 1015
rect 64197 969 64243 1015
rect 64321 969 64367 1015
rect 64445 969 64491 1015
rect 64569 969 64615 1015
rect 64693 969 64739 1015
rect 64817 969 64863 1015
rect 64941 969 64987 1015
rect 65065 969 65111 1015
rect 65189 969 65235 1015
rect 65313 969 65359 1015
rect 65437 969 65483 1015
rect 65561 969 65607 1015
rect 65685 969 65731 1015
rect 65809 969 65855 1015
rect 65933 969 65979 1015
rect 66057 969 66103 1015
rect 66181 969 66227 1015
rect 66305 969 66351 1015
rect 66429 969 66475 1015
rect 66553 969 66599 1015
rect 66677 969 66723 1015
rect 66801 969 66847 1015
rect 66925 969 66971 1015
rect 67049 969 67095 1015
rect 67173 969 67219 1015
rect 67297 969 67343 1015
rect 67421 969 67467 1015
rect 67545 969 67591 1015
rect 67669 969 67715 1015
rect 67793 969 67839 1015
rect 67917 969 67963 1015
rect 68041 969 68087 1015
rect 68165 969 68211 1015
rect 68289 969 68335 1015
rect 68413 969 68459 1015
rect 68537 969 68583 1015
rect 68661 969 68707 1015
rect 68785 969 68831 1015
rect 68909 969 68955 1015
rect 69033 969 69079 1015
rect 69157 969 69203 1015
rect 69281 969 69327 1015
rect 69405 969 69451 1015
rect 69529 969 69575 1015
rect 69653 969 69699 1015
rect 69777 969 69823 1015
rect 69901 969 69947 1015
rect 70025 969 70071 1015
rect 70149 969 70195 1015
rect 70273 969 70319 1015
rect 70397 969 70443 1015
rect 70521 969 70567 1015
rect 70645 969 70691 1015
rect 70769 969 70815 1015
rect 70893 969 70939 1015
rect 71017 969 71063 1015
rect 71141 969 71187 1015
rect 71265 969 71311 1015
rect 71389 969 71435 1015
rect 71513 969 71559 1015
rect 71637 969 71683 1015
rect 71761 969 71807 1015
rect 71885 969 71931 1015
rect 72009 969 72055 1015
rect 72133 969 72179 1015
rect 72257 969 72303 1015
rect 72381 969 72427 1015
rect 72505 969 72551 1015
rect 72629 969 72675 1015
rect 72753 969 72799 1015
rect 72877 969 72923 1015
rect 73001 969 73047 1015
rect 73125 969 73171 1015
rect 73249 969 73295 1015
rect 73373 969 73419 1015
rect 73497 969 73543 1015
rect 73621 969 73667 1015
rect 73745 969 73791 1015
rect 73869 969 73915 1015
rect 73993 969 74039 1015
rect 74117 969 74163 1015
rect 74241 969 74287 1015
rect 74365 969 74411 1015
rect 74489 969 74535 1015
rect 74613 969 74659 1015
rect 74737 969 74783 1015
rect 74861 969 74907 1015
rect 74985 969 75031 1015
rect 75109 969 75155 1015
rect 75233 969 75279 1015
rect 75357 969 75403 1015
rect 75481 969 75527 1015
rect 75605 969 75651 1015
rect 75729 969 75775 1015
rect 75853 969 75899 1015
rect 75977 969 76023 1015
rect 76101 969 76147 1015
rect 76225 969 76271 1015
rect 76349 969 76395 1015
rect 76473 969 76519 1015
rect 76597 969 76643 1015
rect 76721 969 76767 1015
rect 76845 969 76891 1015
rect 76969 969 77015 1015
rect 77093 969 77139 1015
rect 77217 969 77263 1015
rect 77341 969 77387 1015
rect 77465 969 77511 1015
rect 77589 969 77635 1015
rect 77713 969 77759 1015
rect 77837 969 77883 1015
rect 77961 969 78007 1015
rect 78085 969 78131 1015
rect 78209 969 78255 1015
rect 78333 969 78379 1015
rect 78457 969 78503 1015
rect 78581 969 78627 1015
rect 78705 969 78751 1015
rect 78829 969 78875 1015
rect 78953 969 78999 1015
rect 79077 969 79123 1015
rect 79201 969 79247 1015
rect 79325 969 79371 1015
rect 79449 969 79495 1015
rect 79573 969 79619 1015
rect 79697 969 79743 1015
rect 79821 969 79867 1015
rect 79945 969 79991 1015
rect 80069 969 80115 1015
rect 80193 969 80239 1015
rect 80317 969 80363 1015
rect 80441 969 80487 1015
rect 80565 969 80611 1015
rect 80689 969 80735 1015
rect 80813 969 80859 1015
rect 80937 969 80983 1015
rect 81061 969 81107 1015
rect 81185 969 81231 1015
rect 81309 969 81355 1015
rect 81433 969 81479 1015
rect 81557 969 81603 1015
rect 81681 969 81727 1015
rect 81805 969 81851 1015
rect 81929 969 81975 1015
rect 82053 969 82099 1015
rect 82177 969 82223 1015
rect 82301 969 82347 1015
rect 82425 969 82471 1015
rect 82549 969 82595 1015
rect 82673 969 82719 1015
rect 82797 969 82843 1015
rect 82921 969 82967 1015
rect 83045 969 83091 1015
rect 83169 969 83215 1015
rect 83293 969 83339 1015
rect 83417 969 83463 1015
rect 83541 969 83587 1015
rect 83665 969 83711 1015
rect 83789 969 83835 1015
rect 83913 969 83959 1015
rect 84037 969 84083 1015
rect 84161 969 84207 1015
rect 84285 969 84331 1015
rect 84409 969 84455 1015
rect 84533 969 84579 1015
rect 84657 969 84703 1015
rect 84781 969 84827 1015
rect 84905 969 84951 1015
rect 85029 969 85075 1015
rect 85153 969 85199 1015
rect 85277 969 85323 1015
rect 85401 969 85447 1015
rect 85525 969 85571 1015
rect 85649 969 85695 1015
rect 89 845 135 891
rect 213 845 259 891
rect 337 845 383 891
rect 461 845 507 891
rect 585 845 631 891
rect 709 845 755 891
rect 833 845 879 891
rect 957 845 1003 891
rect 1081 845 1127 891
rect 1205 845 1251 891
rect 1329 845 1375 891
rect 1453 845 1499 891
rect 1577 845 1623 891
rect 1701 845 1747 891
rect 1825 845 1871 891
rect 1949 845 1995 891
rect 2073 845 2119 891
rect 2197 845 2243 891
rect 2321 845 2367 891
rect 2445 845 2491 891
rect 2569 845 2615 891
rect 2693 845 2739 891
rect 2817 845 2863 891
rect 2941 845 2987 891
rect 3065 845 3111 891
rect 3189 845 3235 891
rect 3313 845 3359 891
rect 3437 845 3483 891
rect 3561 845 3607 891
rect 3685 845 3731 891
rect 3809 845 3855 891
rect 3933 845 3979 891
rect 4057 845 4103 891
rect 4181 845 4227 891
rect 4305 845 4351 891
rect 4429 845 4475 891
rect 4553 845 4599 891
rect 4677 845 4723 891
rect 4801 845 4847 891
rect 4925 845 4971 891
rect 5049 845 5095 891
rect 5173 845 5219 891
rect 5297 845 5343 891
rect 5421 845 5467 891
rect 5545 845 5591 891
rect 5669 845 5715 891
rect 5793 845 5839 891
rect 5917 845 5963 891
rect 6041 845 6087 891
rect 6165 845 6211 891
rect 6289 845 6335 891
rect 6413 845 6459 891
rect 6537 845 6583 891
rect 6661 845 6707 891
rect 6785 845 6831 891
rect 6909 845 6955 891
rect 7033 845 7079 891
rect 7157 845 7203 891
rect 7281 845 7327 891
rect 7405 845 7451 891
rect 7529 845 7575 891
rect 7653 845 7699 891
rect 7777 845 7823 891
rect 7901 845 7947 891
rect 8025 845 8071 891
rect 8149 845 8195 891
rect 8273 845 8319 891
rect 8397 845 8443 891
rect 8521 845 8567 891
rect 8645 845 8691 891
rect 8769 845 8815 891
rect 8893 845 8939 891
rect 9017 845 9063 891
rect 9141 845 9187 891
rect 9265 845 9311 891
rect 9389 845 9435 891
rect 9513 845 9559 891
rect 9637 845 9683 891
rect 9761 845 9807 891
rect 9885 845 9931 891
rect 10009 845 10055 891
rect 10133 845 10179 891
rect 10257 845 10303 891
rect 10381 845 10427 891
rect 10505 845 10551 891
rect 10629 845 10675 891
rect 10753 845 10799 891
rect 10877 845 10923 891
rect 11001 845 11047 891
rect 11125 845 11171 891
rect 11249 845 11295 891
rect 11373 845 11419 891
rect 11497 845 11543 891
rect 11621 845 11667 891
rect 11745 845 11791 891
rect 11869 845 11915 891
rect 11993 845 12039 891
rect 12117 845 12163 891
rect 12241 845 12287 891
rect 12365 845 12411 891
rect 12489 845 12535 891
rect 12613 845 12659 891
rect 12737 845 12783 891
rect 12861 845 12907 891
rect 12985 845 13031 891
rect 13109 845 13155 891
rect 13233 845 13279 891
rect 13357 845 13403 891
rect 13481 845 13527 891
rect 13605 845 13651 891
rect 13729 845 13775 891
rect 13853 845 13899 891
rect 13977 845 14023 891
rect 14101 845 14147 891
rect 14225 845 14271 891
rect 14349 845 14395 891
rect 14473 845 14519 891
rect 14597 845 14643 891
rect 14721 845 14767 891
rect 14845 845 14891 891
rect 14969 845 15015 891
rect 15093 845 15139 891
rect 15217 845 15263 891
rect 15341 845 15387 891
rect 15465 845 15511 891
rect 15589 845 15635 891
rect 15713 845 15759 891
rect 15837 845 15883 891
rect 15961 845 16007 891
rect 16085 845 16131 891
rect 16209 845 16255 891
rect 16333 845 16379 891
rect 16457 845 16503 891
rect 16581 845 16627 891
rect 16705 845 16751 891
rect 16829 845 16875 891
rect 16953 845 16999 891
rect 17077 845 17123 891
rect 17201 845 17247 891
rect 17325 845 17371 891
rect 17449 845 17495 891
rect 17573 845 17619 891
rect 17697 845 17743 891
rect 17821 845 17867 891
rect 17945 845 17991 891
rect 18069 845 18115 891
rect 18193 845 18239 891
rect 18317 845 18363 891
rect 18441 845 18487 891
rect 18565 845 18611 891
rect 18689 845 18735 891
rect 18813 845 18859 891
rect 18937 845 18983 891
rect 19061 845 19107 891
rect 19185 845 19231 891
rect 19309 845 19355 891
rect 19433 845 19479 891
rect 19557 845 19603 891
rect 19681 845 19727 891
rect 19805 845 19851 891
rect 19929 845 19975 891
rect 20053 845 20099 891
rect 20177 845 20223 891
rect 20301 845 20347 891
rect 20425 845 20471 891
rect 20549 845 20595 891
rect 20673 845 20719 891
rect 20797 845 20843 891
rect 20921 845 20967 891
rect 21045 845 21091 891
rect 21169 845 21215 891
rect 21293 845 21339 891
rect 21417 845 21463 891
rect 21541 845 21587 891
rect 21665 845 21711 891
rect 21789 845 21835 891
rect 21913 845 21959 891
rect 22037 845 22083 891
rect 22161 845 22207 891
rect 22285 845 22331 891
rect 22409 845 22455 891
rect 22533 845 22579 891
rect 22657 845 22703 891
rect 22781 845 22827 891
rect 22905 845 22951 891
rect 23029 845 23075 891
rect 23153 845 23199 891
rect 23277 845 23323 891
rect 23401 845 23447 891
rect 23525 845 23571 891
rect 23649 845 23695 891
rect 23773 845 23819 891
rect 23897 845 23943 891
rect 24021 845 24067 891
rect 24145 845 24191 891
rect 24269 845 24315 891
rect 24393 845 24439 891
rect 24517 845 24563 891
rect 24641 845 24687 891
rect 24765 845 24811 891
rect 24889 845 24935 891
rect 25013 845 25059 891
rect 25137 845 25183 891
rect 25261 845 25307 891
rect 25385 845 25431 891
rect 25509 845 25555 891
rect 25633 845 25679 891
rect 25757 845 25803 891
rect 25881 845 25927 891
rect 26005 845 26051 891
rect 26129 845 26175 891
rect 26253 845 26299 891
rect 26377 845 26423 891
rect 26501 845 26547 891
rect 26625 845 26671 891
rect 26749 845 26795 891
rect 26873 845 26919 891
rect 26997 845 27043 891
rect 27121 845 27167 891
rect 27245 845 27291 891
rect 27369 845 27415 891
rect 27493 845 27539 891
rect 27617 845 27663 891
rect 27741 845 27787 891
rect 27865 845 27911 891
rect 27989 845 28035 891
rect 28113 845 28159 891
rect 28237 845 28283 891
rect 28361 845 28407 891
rect 28485 845 28531 891
rect 28609 845 28655 891
rect 28733 845 28779 891
rect 28857 845 28903 891
rect 28981 845 29027 891
rect 29105 845 29151 891
rect 29229 845 29275 891
rect 29353 845 29399 891
rect 29477 845 29523 891
rect 29601 845 29647 891
rect 29725 845 29771 891
rect 29849 845 29895 891
rect 29973 845 30019 891
rect 30097 845 30143 891
rect 30221 845 30267 891
rect 30345 845 30391 891
rect 30469 845 30515 891
rect 30593 845 30639 891
rect 30717 845 30763 891
rect 30841 845 30887 891
rect 30965 845 31011 891
rect 31089 845 31135 891
rect 31213 845 31259 891
rect 31337 845 31383 891
rect 31461 845 31507 891
rect 31585 845 31631 891
rect 31709 845 31755 891
rect 31833 845 31879 891
rect 31957 845 32003 891
rect 32081 845 32127 891
rect 32205 845 32251 891
rect 32329 845 32375 891
rect 32453 845 32499 891
rect 32577 845 32623 891
rect 32701 845 32747 891
rect 32825 845 32871 891
rect 32949 845 32995 891
rect 33073 845 33119 891
rect 33197 845 33243 891
rect 33321 845 33367 891
rect 33445 845 33491 891
rect 33569 845 33615 891
rect 33693 845 33739 891
rect 33817 845 33863 891
rect 33941 845 33987 891
rect 34065 845 34111 891
rect 34189 845 34235 891
rect 34313 845 34359 891
rect 34437 845 34483 891
rect 34561 845 34607 891
rect 34685 845 34731 891
rect 34809 845 34855 891
rect 34933 845 34979 891
rect 35057 845 35103 891
rect 35181 845 35227 891
rect 35305 845 35351 891
rect 35429 845 35475 891
rect 35553 845 35599 891
rect 35677 845 35723 891
rect 35801 845 35847 891
rect 35925 845 35971 891
rect 36049 845 36095 891
rect 36173 845 36219 891
rect 36297 845 36343 891
rect 36421 845 36467 891
rect 36545 845 36591 891
rect 36669 845 36715 891
rect 36793 845 36839 891
rect 36917 845 36963 891
rect 37041 845 37087 891
rect 37165 845 37211 891
rect 37289 845 37335 891
rect 37413 845 37459 891
rect 37537 845 37583 891
rect 37661 845 37707 891
rect 37785 845 37831 891
rect 37909 845 37955 891
rect 38033 845 38079 891
rect 38157 845 38203 891
rect 38281 845 38327 891
rect 38405 845 38451 891
rect 38529 845 38575 891
rect 38653 845 38699 891
rect 38777 845 38823 891
rect 38901 845 38947 891
rect 39025 845 39071 891
rect 39149 845 39195 891
rect 39273 845 39319 891
rect 39397 845 39443 891
rect 39521 845 39567 891
rect 39645 845 39691 891
rect 39769 845 39815 891
rect 39893 845 39939 891
rect 40017 845 40063 891
rect 40141 845 40187 891
rect 40265 845 40311 891
rect 40389 845 40435 891
rect 40513 845 40559 891
rect 40637 845 40683 891
rect 40761 845 40807 891
rect 40885 845 40931 891
rect 41009 845 41055 891
rect 41133 845 41179 891
rect 41257 845 41303 891
rect 41381 845 41427 891
rect 41505 845 41551 891
rect 41629 845 41675 891
rect 41753 845 41799 891
rect 41877 845 41923 891
rect 42001 845 42047 891
rect 42125 845 42171 891
rect 42249 845 42295 891
rect 42373 845 42419 891
rect 42497 845 42543 891
rect 42621 845 42667 891
rect 42745 845 42791 891
rect 42869 845 42915 891
rect 42993 845 43039 891
rect 43117 845 43163 891
rect 43241 845 43287 891
rect 43365 845 43411 891
rect 43489 845 43535 891
rect 43613 845 43659 891
rect 43737 845 43783 891
rect 43861 845 43907 891
rect 43985 845 44031 891
rect 44109 845 44155 891
rect 44233 845 44279 891
rect 44357 845 44403 891
rect 44481 845 44527 891
rect 44605 845 44651 891
rect 44729 845 44775 891
rect 44853 845 44899 891
rect 44977 845 45023 891
rect 45101 845 45147 891
rect 45225 845 45271 891
rect 45349 845 45395 891
rect 45473 845 45519 891
rect 45597 845 45643 891
rect 45721 845 45767 891
rect 45845 845 45891 891
rect 45969 845 46015 891
rect 46093 845 46139 891
rect 46217 845 46263 891
rect 46341 845 46387 891
rect 46465 845 46511 891
rect 46589 845 46635 891
rect 46713 845 46759 891
rect 46837 845 46883 891
rect 46961 845 47007 891
rect 47085 845 47131 891
rect 47209 845 47255 891
rect 47333 845 47379 891
rect 47457 845 47503 891
rect 47581 845 47627 891
rect 47705 845 47751 891
rect 47829 845 47875 891
rect 47953 845 47999 891
rect 48077 845 48123 891
rect 48201 845 48247 891
rect 48325 845 48371 891
rect 48449 845 48495 891
rect 48573 845 48619 891
rect 48697 845 48743 891
rect 48821 845 48867 891
rect 48945 845 48991 891
rect 49069 845 49115 891
rect 49193 845 49239 891
rect 49317 845 49363 891
rect 49441 845 49487 891
rect 49565 845 49611 891
rect 49689 845 49735 891
rect 49813 845 49859 891
rect 49937 845 49983 891
rect 50061 845 50107 891
rect 50185 845 50231 891
rect 50309 845 50355 891
rect 50433 845 50479 891
rect 50557 845 50603 891
rect 50681 845 50727 891
rect 50805 845 50851 891
rect 50929 845 50975 891
rect 51053 845 51099 891
rect 51177 845 51223 891
rect 51301 845 51347 891
rect 51425 845 51471 891
rect 51549 845 51595 891
rect 51673 845 51719 891
rect 51797 845 51843 891
rect 51921 845 51967 891
rect 52045 845 52091 891
rect 52169 845 52215 891
rect 52293 845 52339 891
rect 52417 845 52463 891
rect 52541 845 52587 891
rect 52665 845 52711 891
rect 52789 845 52835 891
rect 52913 845 52959 891
rect 53037 845 53083 891
rect 53161 845 53207 891
rect 53285 845 53331 891
rect 53409 845 53455 891
rect 53533 845 53579 891
rect 53657 845 53703 891
rect 53781 845 53827 891
rect 53905 845 53951 891
rect 54029 845 54075 891
rect 54153 845 54199 891
rect 54277 845 54323 891
rect 54401 845 54447 891
rect 54525 845 54571 891
rect 54649 845 54695 891
rect 54773 845 54819 891
rect 54897 845 54943 891
rect 55021 845 55067 891
rect 55145 845 55191 891
rect 55269 845 55315 891
rect 55393 845 55439 891
rect 55517 845 55563 891
rect 55641 845 55687 891
rect 55765 845 55811 891
rect 55889 845 55935 891
rect 56013 845 56059 891
rect 56137 845 56183 891
rect 56261 845 56307 891
rect 56385 845 56431 891
rect 56509 845 56555 891
rect 56633 845 56679 891
rect 56757 845 56803 891
rect 56881 845 56927 891
rect 57005 845 57051 891
rect 57129 845 57175 891
rect 57253 845 57299 891
rect 57377 845 57423 891
rect 57501 845 57547 891
rect 57625 845 57671 891
rect 57749 845 57795 891
rect 57873 845 57919 891
rect 57997 845 58043 891
rect 58121 845 58167 891
rect 58245 845 58291 891
rect 58369 845 58415 891
rect 58493 845 58539 891
rect 58617 845 58663 891
rect 58741 845 58787 891
rect 58865 845 58911 891
rect 58989 845 59035 891
rect 59113 845 59159 891
rect 59237 845 59283 891
rect 59361 845 59407 891
rect 59485 845 59531 891
rect 59609 845 59655 891
rect 59733 845 59779 891
rect 59857 845 59903 891
rect 59981 845 60027 891
rect 60105 845 60151 891
rect 60229 845 60275 891
rect 60353 845 60399 891
rect 60477 845 60523 891
rect 60601 845 60647 891
rect 60725 845 60771 891
rect 60849 845 60895 891
rect 60973 845 61019 891
rect 61097 845 61143 891
rect 61221 845 61267 891
rect 61345 845 61391 891
rect 61469 845 61515 891
rect 61593 845 61639 891
rect 61717 845 61763 891
rect 61841 845 61887 891
rect 61965 845 62011 891
rect 62089 845 62135 891
rect 62213 845 62259 891
rect 62337 845 62383 891
rect 62461 845 62507 891
rect 62585 845 62631 891
rect 62709 845 62755 891
rect 62833 845 62879 891
rect 62957 845 63003 891
rect 63081 845 63127 891
rect 63205 845 63251 891
rect 63329 845 63375 891
rect 63453 845 63499 891
rect 63577 845 63623 891
rect 63701 845 63747 891
rect 63825 845 63871 891
rect 63949 845 63995 891
rect 64073 845 64119 891
rect 64197 845 64243 891
rect 64321 845 64367 891
rect 64445 845 64491 891
rect 64569 845 64615 891
rect 64693 845 64739 891
rect 64817 845 64863 891
rect 64941 845 64987 891
rect 65065 845 65111 891
rect 65189 845 65235 891
rect 65313 845 65359 891
rect 65437 845 65483 891
rect 65561 845 65607 891
rect 65685 845 65731 891
rect 65809 845 65855 891
rect 65933 845 65979 891
rect 66057 845 66103 891
rect 66181 845 66227 891
rect 66305 845 66351 891
rect 66429 845 66475 891
rect 66553 845 66599 891
rect 66677 845 66723 891
rect 66801 845 66847 891
rect 66925 845 66971 891
rect 67049 845 67095 891
rect 67173 845 67219 891
rect 67297 845 67343 891
rect 67421 845 67467 891
rect 67545 845 67591 891
rect 67669 845 67715 891
rect 67793 845 67839 891
rect 67917 845 67963 891
rect 68041 845 68087 891
rect 68165 845 68211 891
rect 68289 845 68335 891
rect 68413 845 68459 891
rect 68537 845 68583 891
rect 68661 845 68707 891
rect 68785 845 68831 891
rect 68909 845 68955 891
rect 69033 845 69079 891
rect 69157 845 69203 891
rect 69281 845 69327 891
rect 69405 845 69451 891
rect 69529 845 69575 891
rect 69653 845 69699 891
rect 69777 845 69823 891
rect 69901 845 69947 891
rect 70025 845 70071 891
rect 70149 845 70195 891
rect 70273 845 70319 891
rect 70397 845 70443 891
rect 70521 845 70567 891
rect 70645 845 70691 891
rect 70769 845 70815 891
rect 70893 845 70939 891
rect 71017 845 71063 891
rect 71141 845 71187 891
rect 71265 845 71311 891
rect 71389 845 71435 891
rect 71513 845 71559 891
rect 71637 845 71683 891
rect 71761 845 71807 891
rect 71885 845 71931 891
rect 72009 845 72055 891
rect 72133 845 72179 891
rect 72257 845 72303 891
rect 72381 845 72427 891
rect 72505 845 72551 891
rect 72629 845 72675 891
rect 72753 845 72799 891
rect 72877 845 72923 891
rect 73001 845 73047 891
rect 73125 845 73171 891
rect 73249 845 73295 891
rect 73373 845 73419 891
rect 73497 845 73543 891
rect 73621 845 73667 891
rect 73745 845 73791 891
rect 73869 845 73915 891
rect 73993 845 74039 891
rect 74117 845 74163 891
rect 74241 845 74287 891
rect 74365 845 74411 891
rect 74489 845 74535 891
rect 74613 845 74659 891
rect 74737 845 74783 891
rect 74861 845 74907 891
rect 74985 845 75031 891
rect 75109 845 75155 891
rect 75233 845 75279 891
rect 75357 845 75403 891
rect 75481 845 75527 891
rect 75605 845 75651 891
rect 75729 845 75775 891
rect 75853 845 75899 891
rect 75977 845 76023 891
rect 76101 845 76147 891
rect 76225 845 76271 891
rect 76349 845 76395 891
rect 76473 845 76519 891
rect 76597 845 76643 891
rect 76721 845 76767 891
rect 76845 845 76891 891
rect 76969 845 77015 891
rect 77093 845 77139 891
rect 77217 845 77263 891
rect 77341 845 77387 891
rect 77465 845 77511 891
rect 77589 845 77635 891
rect 77713 845 77759 891
rect 77837 845 77883 891
rect 77961 845 78007 891
rect 78085 845 78131 891
rect 78209 845 78255 891
rect 78333 845 78379 891
rect 78457 845 78503 891
rect 78581 845 78627 891
rect 78705 845 78751 891
rect 78829 845 78875 891
rect 78953 845 78999 891
rect 79077 845 79123 891
rect 79201 845 79247 891
rect 79325 845 79371 891
rect 79449 845 79495 891
rect 79573 845 79619 891
rect 79697 845 79743 891
rect 79821 845 79867 891
rect 79945 845 79991 891
rect 80069 845 80115 891
rect 80193 845 80239 891
rect 80317 845 80363 891
rect 80441 845 80487 891
rect 80565 845 80611 891
rect 80689 845 80735 891
rect 80813 845 80859 891
rect 80937 845 80983 891
rect 81061 845 81107 891
rect 81185 845 81231 891
rect 81309 845 81355 891
rect 81433 845 81479 891
rect 81557 845 81603 891
rect 81681 845 81727 891
rect 81805 845 81851 891
rect 81929 845 81975 891
rect 82053 845 82099 891
rect 82177 845 82223 891
rect 82301 845 82347 891
rect 82425 845 82471 891
rect 82549 845 82595 891
rect 82673 845 82719 891
rect 82797 845 82843 891
rect 82921 845 82967 891
rect 83045 845 83091 891
rect 83169 845 83215 891
rect 83293 845 83339 891
rect 83417 845 83463 891
rect 83541 845 83587 891
rect 83665 845 83711 891
rect 83789 845 83835 891
rect 83913 845 83959 891
rect 84037 845 84083 891
rect 84161 845 84207 891
rect 84285 845 84331 891
rect 84409 845 84455 891
rect 84533 845 84579 891
rect 84657 845 84703 891
rect 84781 845 84827 891
rect 84905 845 84951 891
rect 85029 845 85075 891
rect 85153 845 85199 891
rect 85277 845 85323 891
rect 85401 845 85447 891
rect 85525 845 85571 891
rect 85649 845 85695 891
rect 89 721 135 767
rect 213 721 259 767
rect 337 721 383 767
rect 461 721 507 767
rect 585 721 631 767
rect 709 721 755 767
rect 833 721 879 767
rect 957 721 1003 767
rect 1081 721 1127 767
rect 1205 721 1251 767
rect 1329 721 1375 767
rect 1453 721 1499 767
rect 1577 721 1623 767
rect 1701 721 1747 767
rect 1825 721 1871 767
rect 1949 721 1995 767
rect 2073 721 2119 767
rect 2197 721 2243 767
rect 2321 721 2367 767
rect 2445 721 2491 767
rect 2569 721 2615 767
rect 2693 721 2739 767
rect 2817 721 2863 767
rect 2941 721 2987 767
rect 3065 721 3111 767
rect 3189 721 3235 767
rect 3313 721 3359 767
rect 3437 721 3483 767
rect 3561 721 3607 767
rect 3685 721 3731 767
rect 3809 721 3855 767
rect 3933 721 3979 767
rect 4057 721 4103 767
rect 4181 721 4227 767
rect 4305 721 4351 767
rect 4429 721 4475 767
rect 4553 721 4599 767
rect 4677 721 4723 767
rect 4801 721 4847 767
rect 4925 721 4971 767
rect 5049 721 5095 767
rect 5173 721 5219 767
rect 5297 721 5343 767
rect 5421 721 5467 767
rect 5545 721 5591 767
rect 5669 721 5715 767
rect 5793 721 5839 767
rect 5917 721 5963 767
rect 6041 721 6087 767
rect 6165 721 6211 767
rect 6289 721 6335 767
rect 6413 721 6459 767
rect 6537 721 6583 767
rect 6661 721 6707 767
rect 6785 721 6831 767
rect 6909 721 6955 767
rect 7033 721 7079 767
rect 7157 721 7203 767
rect 7281 721 7327 767
rect 7405 721 7451 767
rect 7529 721 7575 767
rect 7653 721 7699 767
rect 7777 721 7823 767
rect 7901 721 7947 767
rect 8025 721 8071 767
rect 8149 721 8195 767
rect 8273 721 8319 767
rect 8397 721 8443 767
rect 8521 721 8567 767
rect 8645 721 8691 767
rect 8769 721 8815 767
rect 8893 721 8939 767
rect 9017 721 9063 767
rect 9141 721 9187 767
rect 9265 721 9311 767
rect 9389 721 9435 767
rect 9513 721 9559 767
rect 9637 721 9683 767
rect 9761 721 9807 767
rect 9885 721 9931 767
rect 10009 721 10055 767
rect 10133 721 10179 767
rect 10257 721 10303 767
rect 10381 721 10427 767
rect 10505 721 10551 767
rect 10629 721 10675 767
rect 10753 721 10799 767
rect 10877 721 10923 767
rect 11001 721 11047 767
rect 11125 721 11171 767
rect 11249 721 11295 767
rect 11373 721 11419 767
rect 11497 721 11543 767
rect 11621 721 11667 767
rect 11745 721 11791 767
rect 11869 721 11915 767
rect 11993 721 12039 767
rect 12117 721 12163 767
rect 12241 721 12287 767
rect 12365 721 12411 767
rect 12489 721 12535 767
rect 12613 721 12659 767
rect 12737 721 12783 767
rect 12861 721 12907 767
rect 12985 721 13031 767
rect 13109 721 13155 767
rect 13233 721 13279 767
rect 13357 721 13403 767
rect 13481 721 13527 767
rect 13605 721 13651 767
rect 13729 721 13775 767
rect 13853 721 13899 767
rect 13977 721 14023 767
rect 14101 721 14147 767
rect 14225 721 14271 767
rect 14349 721 14395 767
rect 14473 721 14519 767
rect 14597 721 14643 767
rect 14721 721 14767 767
rect 14845 721 14891 767
rect 14969 721 15015 767
rect 15093 721 15139 767
rect 15217 721 15263 767
rect 15341 721 15387 767
rect 15465 721 15511 767
rect 15589 721 15635 767
rect 15713 721 15759 767
rect 15837 721 15883 767
rect 15961 721 16007 767
rect 16085 721 16131 767
rect 16209 721 16255 767
rect 16333 721 16379 767
rect 16457 721 16503 767
rect 16581 721 16627 767
rect 16705 721 16751 767
rect 16829 721 16875 767
rect 16953 721 16999 767
rect 17077 721 17123 767
rect 17201 721 17247 767
rect 17325 721 17371 767
rect 17449 721 17495 767
rect 17573 721 17619 767
rect 17697 721 17743 767
rect 17821 721 17867 767
rect 17945 721 17991 767
rect 18069 721 18115 767
rect 18193 721 18239 767
rect 18317 721 18363 767
rect 18441 721 18487 767
rect 18565 721 18611 767
rect 18689 721 18735 767
rect 18813 721 18859 767
rect 18937 721 18983 767
rect 19061 721 19107 767
rect 19185 721 19231 767
rect 19309 721 19355 767
rect 19433 721 19479 767
rect 19557 721 19603 767
rect 19681 721 19727 767
rect 19805 721 19851 767
rect 19929 721 19975 767
rect 20053 721 20099 767
rect 20177 721 20223 767
rect 20301 721 20347 767
rect 20425 721 20471 767
rect 20549 721 20595 767
rect 20673 721 20719 767
rect 20797 721 20843 767
rect 20921 721 20967 767
rect 21045 721 21091 767
rect 21169 721 21215 767
rect 21293 721 21339 767
rect 21417 721 21463 767
rect 21541 721 21587 767
rect 21665 721 21711 767
rect 21789 721 21835 767
rect 21913 721 21959 767
rect 22037 721 22083 767
rect 22161 721 22207 767
rect 22285 721 22331 767
rect 22409 721 22455 767
rect 22533 721 22579 767
rect 22657 721 22703 767
rect 22781 721 22827 767
rect 22905 721 22951 767
rect 23029 721 23075 767
rect 23153 721 23199 767
rect 23277 721 23323 767
rect 23401 721 23447 767
rect 23525 721 23571 767
rect 23649 721 23695 767
rect 23773 721 23819 767
rect 23897 721 23943 767
rect 24021 721 24067 767
rect 24145 721 24191 767
rect 24269 721 24315 767
rect 24393 721 24439 767
rect 24517 721 24563 767
rect 24641 721 24687 767
rect 24765 721 24811 767
rect 24889 721 24935 767
rect 25013 721 25059 767
rect 25137 721 25183 767
rect 25261 721 25307 767
rect 25385 721 25431 767
rect 25509 721 25555 767
rect 25633 721 25679 767
rect 25757 721 25803 767
rect 25881 721 25927 767
rect 26005 721 26051 767
rect 26129 721 26175 767
rect 26253 721 26299 767
rect 26377 721 26423 767
rect 26501 721 26547 767
rect 26625 721 26671 767
rect 26749 721 26795 767
rect 26873 721 26919 767
rect 26997 721 27043 767
rect 27121 721 27167 767
rect 27245 721 27291 767
rect 27369 721 27415 767
rect 27493 721 27539 767
rect 27617 721 27663 767
rect 27741 721 27787 767
rect 27865 721 27911 767
rect 27989 721 28035 767
rect 28113 721 28159 767
rect 28237 721 28283 767
rect 28361 721 28407 767
rect 28485 721 28531 767
rect 28609 721 28655 767
rect 28733 721 28779 767
rect 28857 721 28903 767
rect 28981 721 29027 767
rect 29105 721 29151 767
rect 29229 721 29275 767
rect 29353 721 29399 767
rect 29477 721 29523 767
rect 29601 721 29647 767
rect 29725 721 29771 767
rect 29849 721 29895 767
rect 29973 721 30019 767
rect 30097 721 30143 767
rect 30221 721 30267 767
rect 30345 721 30391 767
rect 30469 721 30515 767
rect 30593 721 30639 767
rect 30717 721 30763 767
rect 30841 721 30887 767
rect 30965 721 31011 767
rect 31089 721 31135 767
rect 31213 721 31259 767
rect 31337 721 31383 767
rect 31461 721 31507 767
rect 31585 721 31631 767
rect 31709 721 31755 767
rect 31833 721 31879 767
rect 31957 721 32003 767
rect 32081 721 32127 767
rect 32205 721 32251 767
rect 32329 721 32375 767
rect 32453 721 32499 767
rect 32577 721 32623 767
rect 32701 721 32747 767
rect 32825 721 32871 767
rect 32949 721 32995 767
rect 33073 721 33119 767
rect 33197 721 33243 767
rect 33321 721 33367 767
rect 33445 721 33491 767
rect 33569 721 33615 767
rect 33693 721 33739 767
rect 33817 721 33863 767
rect 33941 721 33987 767
rect 34065 721 34111 767
rect 34189 721 34235 767
rect 34313 721 34359 767
rect 34437 721 34483 767
rect 34561 721 34607 767
rect 34685 721 34731 767
rect 34809 721 34855 767
rect 34933 721 34979 767
rect 35057 721 35103 767
rect 35181 721 35227 767
rect 35305 721 35351 767
rect 35429 721 35475 767
rect 35553 721 35599 767
rect 35677 721 35723 767
rect 35801 721 35847 767
rect 35925 721 35971 767
rect 36049 721 36095 767
rect 36173 721 36219 767
rect 36297 721 36343 767
rect 36421 721 36467 767
rect 36545 721 36591 767
rect 36669 721 36715 767
rect 36793 721 36839 767
rect 36917 721 36963 767
rect 37041 721 37087 767
rect 37165 721 37211 767
rect 37289 721 37335 767
rect 37413 721 37459 767
rect 37537 721 37583 767
rect 37661 721 37707 767
rect 37785 721 37831 767
rect 37909 721 37955 767
rect 38033 721 38079 767
rect 38157 721 38203 767
rect 38281 721 38327 767
rect 38405 721 38451 767
rect 38529 721 38575 767
rect 38653 721 38699 767
rect 38777 721 38823 767
rect 38901 721 38947 767
rect 39025 721 39071 767
rect 39149 721 39195 767
rect 39273 721 39319 767
rect 39397 721 39443 767
rect 39521 721 39567 767
rect 39645 721 39691 767
rect 39769 721 39815 767
rect 39893 721 39939 767
rect 40017 721 40063 767
rect 40141 721 40187 767
rect 40265 721 40311 767
rect 40389 721 40435 767
rect 40513 721 40559 767
rect 40637 721 40683 767
rect 40761 721 40807 767
rect 40885 721 40931 767
rect 41009 721 41055 767
rect 41133 721 41179 767
rect 41257 721 41303 767
rect 41381 721 41427 767
rect 41505 721 41551 767
rect 41629 721 41675 767
rect 41753 721 41799 767
rect 41877 721 41923 767
rect 42001 721 42047 767
rect 42125 721 42171 767
rect 42249 721 42295 767
rect 42373 721 42419 767
rect 42497 721 42543 767
rect 42621 721 42667 767
rect 42745 721 42791 767
rect 42869 721 42915 767
rect 42993 721 43039 767
rect 43117 721 43163 767
rect 43241 721 43287 767
rect 43365 721 43411 767
rect 43489 721 43535 767
rect 43613 721 43659 767
rect 43737 721 43783 767
rect 43861 721 43907 767
rect 43985 721 44031 767
rect 44109 721 44155 767
rect 44233 721 44279 767
rect 44357 721 44403 767
rect 44481 721 44527 767
rect 44605 721 44651 767
rect 44729 721 44775 767
rect 44853 721 44899 767
rect 44977 721 45023 767
rect 45101 721 45147 767
rect 45225 721 45271 767
rect 45349 721 45395 767
rect 45473 721 45519 767
rect 45597 721 45643 767
rect 45721 721 45767 767
rect 45845 721 45891 767
rect 45969 721 46015 767
rect 46093 721 46139 767
rect 46217 721 46263 767
rect 46341 721 46387 767
rect 46465 721 46511 767
rect 46589 721 46635 767
rect 46713 721 46759 767
rect 46837 721 46883 767
rect 46961 721 47007 767
rect 47085 721 47131 767
rect 47209 721 47255 767
rect 47333 721 47379 767
rect 47457 721 47503 767
rect 47581 721 47627 767
rect 47705 721 47751 767
rect 47829 721 47875 767
rect 47953 721 47999 767
rect 48077 721 48123 767
rect 48201 721 48247 767
rect 48325 721 48371 767
rect 48449 721 48495 767
rect 48573 721 48619 767
rect 48697 721 48743 767
rect 48821 721 48867 767
rect 48945 721 48991 767
rect 49069 721 49115 767
rect 49193 721 49239 767
rect 49317 721 49363 767
rect 49441 721 49487 767
rect 49565 721 49611 767
rect 49689 721 49735 767
rect 49813 721 49859 767
rect 49937 721 49983 767
rect 50061 721 50107 767
rect 50185 721 50231 767
rect 50309 721 50355 767
rect 50433 721 50479 767
rect 50557 721 50603 767
rect 50681 721 50727 767
rect 50805 721 50851 767
rect 50929 721 50975 767
rect 51053 721 51099 767
rect 51177 721 51223 767
rect 51301 721 51347 767
rect 51425 721 51471 767
rect 51549 721 51595 767
rect 51673 721 51719 767
rect 51797 721 51843 767
rect 51921 721 51967 767
rect 52045 721 52091 767
rect 52169 721 52215 767
rect 52293 721 52339 767
rect 52417 721 52463 767
rect 52541 721 52587 767
rect 52665 721 52711 767
rect 52789 721 52835 767
rect 52913 721 52959 767
rect 53037 721 53083 767
rect 53161 721 53207 767
rect 53285 721 53331 767
rect 53409 721 53455 767
rect 53533 721 53579 767
rect 53657 721 53703 767
rect 53781 721 53827 767
rect 53905 721 53951 767
rect 54029 721 54075 767
rect 54153 721 54199 767
rect 54277 721 54323 767
rect 54401 721 54447 767
rect 54525 721 54571 767
rect 54649 721 54695 767
rect 54773 721 54819 767
rect 54897 721 54943 767
rect 55021 721 55067 767
rect 55145 721 55191 767
rect 55269 721 55315 767
rect 55393 721 55439 767
rect 55517 721 55563 767
rect 55641 721 55687 767
rect 55765 721 55811 767
rect 55889 721 55935 767
rect 56013 721 56059 767
rect 56137 721 56183 767
rect 56261 721 56307 767
rect 56385 721 56431 767
rect 56509 721 56555 767
rect 56633 721 56679 767
rect 56757 721 56803 767
rect 56881 721 56927 767
rect 57005 721 57051 767
rect 57129 721 57175 767
rect 57253 721 57299 767
rect 57377 721 57423 767
rect 57501 721 57547 767
rect 57625 721 57671 767
rect 57749 721 57795 767
rect 57873 721 57919 767
rect 57997 721 58043 767
rect 58121 721 58167 767
rect 58245 721 58291 767
rect 58369 721 58415 767
rect 58493 721 58539 767
rect 58617 721 58663 767
rect 58741 721 58787 767
rect 58865 721 58911 767
rect 58989 721 59035 767
rect 59113 721 59159 767
rect 59237 721 59283 767
rect 59361 721 59407 767
rect 59485 721 59531 767
rect 59609 721 59655 767
rect 59733 721 59779 767
rect 59857 721 59903 767
rect 59981 721 60027 767
rect 60105 721 60151 767
rect 60229 721 60275 767
rect 60353 721 60399 767
rect 60477 721 60523 767
rect 60601 721 60647 767
rect 60725 721 60771 767
rect 60849 721 60895 767
rect 60973 721 61019 767
rect 61097 721 61143 767
rect 61221 721 61267 767
rect 61345 721 61391 767
rect 61469 721 61515 767
rect 61593 721 61639 767
rect 61717 721 61763 767
rect 61841 721 61887 767
rect 61965 721 62011 767
rect 62089 721 62135 767
rect 62213 721 62259 767
rect 62337 721 62383 767
rect 62461 721 62507 767
rect 62585 721 62631 767
rect 62709 721 62755 767
rect 62833 721 62879 767
rect 62957 721 63003 767
rect 63081 721 63127 767
rect 63205 721 63251 767
rect 63329 721 63375 767
rect 63453 721 63499 767
rect 63577 721 63623 767
rect 63701 721 63747 767
rect 63825 721 63871 767
rect 63949 721 63995 767
rect 64073 721 64119 767
rect 64197 721 64243 767
rect 64321 721 64367 767
rect 64445 721 64491 767
rect 64569 721 64615 767
rect 64693 721 64739 767
rect 64817 721 64863 767
rect 64941 721 64987 767
rect 65065 721 65111 767
rect 65189 721 65235 767
rect 65313 721 65359 767
rect 65437 721 65483 767
rect 65561 721 65607 767
rect 65685 721 65731 767
rect 65809 721 65855 767
rect 65933 721 65979 767
rect 66057 721 66103 767
rect 66181 721 66227 767
rect 66305 721 66351 767
rect 66429 721 66475 767
rect 66553 721 66599 767
rect 66677 721 66723 767
rect 66801 721 66847 767
rect 66925 721 66971 767
rect 67049 721 67095 767
rect 67173 721 67219 767
rect 67297 721 67343 767
rect 67421 721 67467 767
rect 67545 721 67591 767
rect 67669 721 67715 767
rect 67793 721 67839 767
rect 67917 721 67963 767
rect 68041 721 68087 767
rect 68165 721 68211 767
rect 68289 721 68335 767
rect 68413 721 68459 767
rect 68537 721 68583 767
rect 68661 721 68707 767
rect 68785 721 68831 767
rect 68909 721 68955 767
rect 69033 721 69079 767
rect 69157 721 69203 767
rect 69281 721 69327 767
rect 69405 721 69451 767
rect 69529 721 69575 767
rect 69653 721 69699 767
rect 69777 721 69823 767
rect 69901 721 69947 767
rect 70025 721 70071 767
rect 70149 721 70195 767
rect 70273 721 70319 767
rect 70397 721 70443 767
rect 70521 721 70567 767
rect 70645 721 70691 767
rect 70769 721 70815 767
rect 70893 721 70939 767
rect 71017 721 71063 767
rect 71141 721 71187 767
rect 71265 721 71311 767
rect 71389 721 71435 767
rect 71513 721 71559 767
rect 71637 721 71683 767
rect 71761 721 71807 767
rect 71885 721 71931 767
rect 72009 721 72055 767
rect 72133 721 72179 767
rect 72257 721 72303 767
rect 72381 721 72427 767
rect 72505 721 72551 767
rect 72629 721 72675 767
rect 72753 721 72799 767
rect 72877 721 72923 767
rect 73001 721 73047 767
rect 73125 721 73171 767
rect 73249 721 73295 767
rect 73373 721 73419 767
rect 73497 721 73543 767
rect 73621 721 73667 767
rect 73745 721 73791 767
rect 73869 721 73915 767
rect 73993 721 74039 767
rect 74117 721 74163 767
rect 74241 721 74287 767
rect 74365 721 74411 767
rect 74489 721 74535 767
rect 74613 721 74659 767
rect 74737 721 74783 767
rect 74861 721 74907 767
rect 74985 721 75031 767
rect 75109 721 75155 767
rect 75233 721 75279 767
rect 75357 721 75403 767
rect 75481 721 75527 767
rect 75605 721 75651 767
rect 75729 721 75775 767
rect 75853 721 75899 767
rect 75977 721 76023 767
rect 76101 721 76147 767
rect 76225 721 76271 767
rect 76349 721 76395 767
rect 76473 721 76519 767
rect 76597 721 76643 767
rect 76721 721 76767 767
rect 76845 721 76891 767
rect 76969 721 77015 767
rect 77093 721 77139 767
rect 77217 721 77263 767
rect 77341 721 77387 767
rect 77465 721 77511 767
rect 77589 721 77635 767
rect 77713 721 77759 767
rect 77837 721 77883 767
rect 77961 721 78007 767
rect 78085 721 78131 767
rect 78209 721 78255 767
rect 78333 721 78379 767
rect 78457 721 78503 767
rect 78581 721 78627 767
rect 78705 721 78751 767
rect 78829 721 78875 767
rect 78953 721 78999 767
rect 79077 721 79123 767
rect 79201 721 79247 767
rect 79325 721 79371 767
rect 79449 721 79495 767
rect 79573 721 79619 767
rect 79697 721 79743 767
rect 79821 721 79867 767
rect 79945 721 79991 767
rect 80069 721 80115 767
rect 80193 721 80239 767
rect 80317 721 80363 767
rect 80441 721 80487 767
rect 80565 721 80611 767
rect 80689 721 80735 767
rect 80813 721 80859 767
rect 80937 721 80983 767
rect 81061 721 81107 767
rect 81185 721 81231 767
rect 81309 721 81355 767
rect 81433 721 81479 767
rect 81557 721 81603 767
rect 81681 721 81727 767
rect 81805 721 81851 767
rect 81929 721 81975 767
rect 82053 721 82099 767
rect 82177 721 82223 767
rect 82301 721 82347 767
rect 82425 721 82471 767
rect 82549 721 82595 767
rect 82673 721 82719 767
rect 82797 721 82843 767
rect 82921 721 82967 767
rect 83045 721 83091 767
rect 83169 721 83215 767
rect 83293 721 83339 767
rect 83417 721 83463 767
rect 83541 721 83587 767
rect 83665 721 83711 767
rect 83789 721 83835 767
rect 83913 721 83959 767
rect 84037 721 84083 767
rect 84161 721 84207 767
rect 84285 721 84331 767
rect 84409 721 84455 767
rect 84533 721 84579 767
rect 84657 721 84703 767
rect 84781 721 84827 767
rect 84905 721 84951 767
rect 85029 721 85075 767
rect 85153 721 85199 767
rect 85277 721 85323 767
rect 85401 721 85447 767
rect 85525 721 85571 767
rect 85649 721 85695 767
rect 89 597 135 643
rect 213 597 259 643
rect 337 597 383 643
rect 461 597 507 643
rect 585 597 631 643
rect 709 597 755 643
rect 833 597 879 643
rect 957 597 1003 643
rect 1081 597 1127 643
rect 1205 597 1251 643
rect 1329 597 1375 643
rect 1453 597 1499 643
rect 1577 597 1623 643
rect 1701 597 1747 643
rect 1825 597 1871 643
rect 1949 597 1995 643
rect 2073 597 2119 643
rect 2197 597 2243 643
rect 2321 597 2367 643
rect 2445 597 2491 643
rect 2569 597 2615 643
rect 2693 597 2739 643
rect 2817 597 2863 643
rect 2941 597 2987 643
rect 3065 597 3111 643
rect 3189 597 3235 643
rect 3313 597 3359 643
rect 3437 597 3483 643
rect 3561 597 3607 643
rect 3685 597 3731 643
rect 3809 597 3855 643
rect 3933 597 3979 643
rect 4057 597 4103 643
rect 4181 597 4227 643
rect 4305 597 4351 643
rect 4429 597 4475 643
rect 4553 597 4599 643
rect 4677 597 4723 643
rect 4801 597 4847 643
rect 4925 597 4971 643
rect 5049 597 5095 643
rect 5173 597 5219 643
rect 5297 597 5343 643
rect 5421 597 5467 643
rect 5545 597 5591 643
rect 5669 597 5715 643
rect 5793 597 5839 643
rect 5917 597 5963 643
rect 6041 597 6087 643
rect 6165 597 6211 643
rect 6289 597 6335 643
rect 6413 597 6459 643
rect 6537 597 6583 643
rect 6661 597 6707 643
rect 6785 597 6831 643
rect 6909 597 6955 643
rect 7033 597 7079 643
rect 7157 597 7203 643
rect 7281 597 7327 643
rect 7405 597 7451 643
rect 7529 597 7575 643
rect 7653 597 7699 643
rect 7777 597 7823 643
rect 7901 597 7947 643
rect 8025 597 8071 643
rect 8149 597 8195 643
rect 8273 597 8319 643
rect 8397 597 8443 643
rect 8521 597 8567 643
rect 8645 597 8691 643
rect 8769 597 8815 643
rect 8893 597 8939 643
rect 9017 597 9063 643
rect 9141 597 9187 643
rect 9265 597 9311 643
rect 9389 597 9435 643
rect 9513 597 9559 643
rect 9637 597 9683 643
rect 9761 597 9807 643
rect 9885 597 9931 643
rect 10009 597 10055 643
rect 10133 597 10179 643
rect 10257 597 10303 643
rect 10381 597 10427 643
rect 10505 597 10551 643
rect 10629 597 10675 643
rect 10753 597 10799 643
rect 10877 597 10923 643
rect 11001 597 11047 643
rect 11125 597 11171 643
rect 11249 597 11295 643
rect 11373 597 11419 643
rect 11497 597 11543 643
rect 11621 597 11667 643
rect 11745 597 11791 643
rect 11869 597 11915 643
rect 11993 597 12039 643
rect 12117 597 12163 643
rect 12241 597 12287 643
rect 12365 597 12411 643
rect 12489 597 12535 643
rect 12613 597 12659 643
rect 12737 597 12783 643
rect 12861 597 12907 643
rect 12985 597 13031 643
rect 13109 597 13155 643
rect 13233 597 13279 643
rect 13357 597 13403 643
rect 13481 597 13527 643
rect 13605 597 13651 643
rect 13729 597 13775 643
rect 13853 597 13899 643
rect 13977 597 14023 643
rect 14101 597 14147 643
rect 14225 597 14271 643
rect 14349 597 14395 643
rect 14473 597 14519 643
rect 14597 597 14643 643
rect 14721 597 14767 643
rect 14845 597 14891 643
rect 14969 597 15015 643
rect 15093 597 15139 643
rect 15217 597 15263 643
rect 15341 597 15387 643
rect 15465 597 15511 643
rect 15589 597 15635 643
rect 15713 597 15759 643
rect 15837 597 15883 643
rect 15961 597 16007 643
rect 16085 597 16131 643
rect 16209 597 16255 643
rect 16333 597 16379 643
rect 16457 597 16503 643
rect 16581 597 16627 643
rect 16705 597 16751 643
rect 16829 597 16875 643
rect 16953 597 16999 643
rect 17077 597 17123 643
rect 17201 597 17247 643
rect 17325 597 17371 643
rect 17449 597 17495 643
rect 17573 597 17619 643
rect 17697 597 17743 643
rect 17821 597 17867 643
rect 17945 597 17991 643
rect 18069 597 18115 643
rect 18193 597 18239 643
rect 18317 597 18363 643
rect 18441 597 18487 643
rect 18565 597 18611 643
rect 18689 597 18735 643
rect 18813 597 18859 643
rect 18937 597 18983 643
rect 19061 597 19107 643
rect 19185 597 19231 643
rect 19309 597 19355 643
rect 19433 597 19479 643
rect 19557 597 19603 643
rect 19681 597 19727 643
rect 19805 597 19851 643
rect 19929 597 19975 643
rect 20053 597 20099 643
rect 20177 597 20223 643
rect 20301 597 20347 643
rect 20425 597 20471 643
rect 20549 597 20595 643
rect 20673 597 20719 643
rect 20797 597 20843 643
rect 20921 597 20967 643
rect 21045 597 21091 643
rect 21169 597 21215 643
rect 21293 597 21339 643
rect 21417 597 21463 643
rect 21541 597 21587 643
rect 21665 597 21711 643
rect 21789 597 21835 643
rect 21913 597 21959 643
rect 22037 597 22083 643
rect 22161 597 22207 643
rect 22285 597 22331 643
rect 22409 597 22455 643
rect 22533 597 22579 643
rect 22657 597 22703 643
rect 22781 597 22827 643
rect 22905 597 22951 643
rect 23029 597 23075 643
rect 23153 597 23199 643
rect 23277 597 23323 643
rect 23401 597 23447 643
rect 23525 597 23571 643
rect 23649 597 23695 643
rect 23773 597 23819 643
rect 23897 597 23943 643
rect 24021 597 24067 643
rect 24145 597 24191 643
rect 24269 597 24315 643
rect 24393 597 24439 643
rect 24517 597 24563 643
rect 24641 597 24687 643
rect 24765 597 24811 643
rect 24889 597 24935 643
rect 25013 597 25059 643
rect 25137 597 25183 643
rect 25261 597 25307 643
rect 25385 597 25431 643
rect 25509 597 25555 643
rect 25633 597 25679 643
rect 25757 597 25803 643
rect 25881 597 25927 643
rect 26005 597 26051 643
rect 26129 597 26175 643
rect 26253 597 26299 643
rect 26377 597 26423 643
rect 26501 597 26547 643
rect 26625 597 26671 643
rect 26749 597 26795 643
rect 26873 597 26919 643
rect 26997 597 27043 643
rect 27121 597 27167 643
rect 27245 597 27291 643
rect 27369 597 27415 643
rect 27493 597 27539 643
rect 27617 597 27663 643
rect 27741 597 27787 643
rect 27865 597 27911 643
rect 27989 597 28035 643
rect 28113 597 28159 643
rect 28237 597 28283 643
rect 28361 597 28407 643
rect 28485 597 28531 643
rect 28609 597 28655 643
rect 28733 597 28779 643
rect 28857 597 28903 643
rect 28981 597 29027 643
rect 29105 597 29151 643
rect 29229 597 29275 643
rect 29353 597 29399 643
rect 29477 597 29523 643
rect 29601 597 29647 643
rect 29725 597 29771 643
rect 29849 597 29895 643
rect 29973 597 30019 643
rect 30097 597 30143 643
rect 30221 597 30267 643
rect 30345 597 30391 643
rect 30469 597 30515 643
rect 30593 597 30639 643
rect 30717 597 30763 643
rect 30841 597 30887 643
rect 30965 597 31011 643
rect 31089 597 31135 643
rect 31213 597 31259 643
rect 31337 597 31383 643
rect 31461 597 31507 643
rect 31585 597 31631 643
rect 31709 597 31755 643
rect 31833 597 31879 643
rect 31957 597 32003 643
rect 32081 597 32127 643
rect 32205 597 32251 643
rect 32329 597 32375 643
rect 32453 597 32499 643
rect 32577 597 32623 643
rect 32701 597 32747 643
rect 32825 597 32871 643
rect 32949 597 32995 643
rect 33073 597 33119 643
rect 33197 597 33243 643
rect 33321 597 33367 643
rect 33445 597 33491 643
rect 33569 597 33615 643
rect 33693 597 33739 643
rect 33817 597 33863 643
rect 33941 597 33987 643
rect 34065 597 34111 643
rect 34189 597 34235 643
rect 34313 597 34359 643
rect 34437 597 34483 643
rect 34561 597 34607 643
rect 34685 597 34731 643
rect 34809 597 34855 643
rect 34933 597 34979 643
rect 35057 597 35103 643
rect 35181 597 35227 643
rect 35305 597 35351 643
rect 35429 597 35475 643
rect 35553 597 35599 643
rect 35677 597 35723 643
rect 35801 597 35847 643
rect 35925 597 35971 643
rect 36049 597 36095 643
rect 36173 597 36219 643
rect 36297 597 36343 643
rect 36421 597 36467 643
rect 36545 597 36591 643
rect 36669 597 36715 643
rect 36793 597 36839 643
rect 36917 597 36963 643
rect 37041 597 37087 643
rect 37165 597 37211 643
rect 37289 597 37335 643
rect 37413 597 37459 643
rect 37537 597 37583 643
rect 37661 597 37707 643
rect 37785 597 37831 643
rect 37909 597 37955 643
rect 38033 597 38079 643
rect 38157 597 38203 643
rect 38281 597 38327 643
rect 38405 597 38451 643
rect 38529 597 38575 643
rect 38653 597 38699 643
rect 38777 597 38823 643
rect 38901 597 38947 643
rect 39025 597 39071 643
rect 39149 597 39195 643
rect 39273 597 39319 643
rect 39397 597 39443 643
rect 39521 597 39567 643
rect 39645 597 39691 643
rect 39769 597 39815 643
rect 39893 597 39939 643
rect 40017 597 40063 643
rect 40141 597 40187 643
rect 40265 597 40311 643
rect 40389 597 40435 643
rect 40513 597 40559 643
rect 40637 597 40683 643
rect 40761 597 40807 643
rect 40885 597 40931 643
rect 41009 597 41055 643
rect 41133 597 41179 643
rect 41257 597 41303 643
rect 41381 597 41427 643
rect 41505 597 41551 643
rect 41629 597 41675 643
rect 41753 597 41799 643
rect 41877 597 41923 643
rect 42001 597 42047 643
rect 42125 597 42171 643
rect 42249 597 42295 643
rect 42373 597 42419 643
rect 42497 597 42543 643
rect 42621 597 42667 643
rect 42745 597 42791 643
rect 42869 597 42915 643
rect 42993 597 43039 643
rect 43117 597 43163 643
rect 43241 597 43287 643
rect 43365 597 43411 643
rect 43489 597 43535 643
rect 43613 597 43659 643
rect 43737 597 43783 643
rect 43861 597 43907 643
rect 43985 597 44031 643
rect 44109 597 44155 643
rect 44233 597 44279 643
rect 44357 597 44403 643
rect 44481 597 44527 643
rect 44605 597 44651 643
rect 44729 597 44775 643
rect 44853 597 44899 643
rect 44977 597 45023 643
rect 45101 597 45147 643
rect 45225 597 45271 643
rect 45349 597 45395 643
rect 45473 597 45519 643
rect 45597 597 45643 643
rect 45721 597 45767 643
rect 45845 597 45891 643
rect 45969 597 46015 643
rect 46093 597 46139 643
rect 46217 597 46263 643
rect 46341 597 46387 643
rect 46465 597 46511 643
rect 46589 597 46635 643
rect 46713 597 46759 643
rect 46837 597 46883 643
rect 46961 597 47007 643
rect 47085 597 47131 643
rect 47209 597 47255 643
rect 47333 597 47379 643
rect 47457 597 47503 643
rect 47581 597 47627 643
rect 47705 597 47751 643
rect 47829 597 47875 643
rect 47953 597 47999 643
rect 48077 597 48123 643
rect 48201 597 48247 643
rect 48325 597 48371 643
rect 48449 597 48495 643
rect 48573 597 48619 643
rect 48697 597 48743 643
rect 48821 597 48867 643
rect 48945 597 48991 643
rect 49069 597 49115 643
rect 49193 597 49239 643
rect 49317 597 49363 643
rect 49441 597 49487 643
rect 49565 597 49611 643
rect 49689 597 49735 643
rect 49813 597 49859 643
rect 49937 597 49983 643
rect 50061 597 50107 643
rect 50185 597 50231 643
rect 50309 597 50355 643
rect 50433 597 50479 643
rect 50557 597 50603 643
rect 50681 597 50727 643
rect 50805 597 50851 643
rect 50929 597 50975 643
rect 51053 597 51099 643
rect 51177 597 51223 643
rect 51301 597 51347 643
rect 51425 597 51471 643
rect 51549 597 51595 643
rect 51673 597 51719 643
rect 51797 597 51843 643
rect 51921 597 51967 643
rect 52045 597 52091 643
rect 52169 597 52215 643
rect 52293 597 52339 643
rect 52417 597 52463 643
rect 52541 597 52587 643
rect 52665 597 52711 643
rect 52789 597 52835 643
rect 52913 597 52959 643
rect 53037 597 53083 643
rect 53161 597 53207 643
rect 53285 597 53331 643
rect 53409 597 53455 643
rect 53533 597 53579 643
rect 53657 597 53703 643
rect 53781 597 53827 643
rect 53905 597 53951 643
rect 54029 597 54075 643
rect 54153 597 54199 643
rect 54277 597 54323 643
rect 54401 597 54447 643
rect 54525 597 54571 643
rect 54649 597 54695 643
rect 54773 597 54819 643
rect 54897 597 54943 643
rect 55021 597 55067 643
rect 55145 597 55191 643
rect 55269 597 55315 643
rect 55393 597 55439 643
rect 55517 597 55563 643
rect 55641 597 55687 643
rect 55765 597 55811 643
rect 55889 597 55935 643
rect 56013 597 56059 643
rect 56137 597 56183 643
rect 56261 597 56307 643
rect 56385 597 56431 643
rect 56509 597 56555 643
rect 56633 597 56679 643
rect 56757 597 56803 643
rect 56881 597 56927 643
rect 57005 597 57051 643
rect 57129 597 57175 643
rect 57253 597 57299 643
rect 57377 597 57423 643
rect 57501 597 57547 643
rect 57625 597 57671 643
rect 57749 597 57795 643
rect 57873 597 57919 643
rect 57997 597 58043 643
rect 58121 597 58167 643
rect 58245 597 58291 643
rect 58369 597 58415 643
rect 58493 597 58539 643
rect 58617 597 58663 643
rect 58741 597 58787 643
rect 58865 597 58911 643
rect 58989 597 59035 643
rect 59113 597 59159 643
rect 59237 597 59283 643
rect 59361 597 59407 643
rect 59485 597 59531 643
rect 59609 597 59655 643
rect 59733 597 59779 643
rect 59857 597 59903 643
rect 59981 597 60027 643
rect 60105 597 60151 643
rect 60229 597 60275 643
rect 60353 597 60399 643
rect 60477 597 60523 643
rect 60601 597 60647 643
rect 60725 597 60771 643
rect 60849 597 60895 643
rect 60973 597 61019 643
rect 61097 597 61143 643
rect 61221 597 61267 643
rect 61345 597 61391 643
rect 61469 597 61515 643
rect 61593 597 61639 643
rect 61717 597 61763 643
rect 61841 597 61887 643
rect 61965 597 62011 643
rect 62089 597 62135 643
rect 62213 597 62259 643
rect 62337 597 62383 643
rect 62461 597 62507 643
rect 62585 597 62631 643
rect 62709 597 62755 643
rect 62833 597 62879 643
rect 62957 597 63003 643
rect 63081 597 63127 643
rect 63205 597 63251 643
rect 63329 597 63375 643
rect 63453 597 63499 643
rect 63577 597 63623 643
rect 63701 597 63747 643
rect 63825 597 63871 643
rect 63949 597 63995 643
rect 64073 597 64119 643
rect 64197 597 64243 643
rect 64321 597 64367 643
rect 64445 597 64491 643
rect 64569 597 64615 643
rect 64693 597 64739 643
rect 64817 597 64863 643
rect 64941 597 64987 643
rect 65065 597 65111 643
rect 65189 597 65235 643
rect 65313 597 65359 643
rect 65437 597 65483 643
rect 65561 597 65607 643
rect 65685 597 65731 643
rect 65809 597 65855 643
rect 65933 597 65979 643
rect 66057 597 66103 643
rect 66181 597 66227 643
rect 66305 597 66351 643
rect 66429 597 66475 643
rect 66553 597 66599 643
rect 66677 597 66723 643
rect 66801 597 66847 643
rect 66925 597 66971 643
rect 67049 597 67095 643
rect 67173 597 67219 643
rect 67297 597 67343 643
rect 67421 597 67467 643
rect 67545 597 67591 643
rect 67669 597 67715 643
rect 67793 597 67839 643
rect 67917 597 67963 643
rect 68041 597 68087 643
rect 68165 597 68211 643
rect 68289 597 68335 643
rect 68413 597 68459 643
rect 68537 597 68583 643
rect 68661 597 68707 643
rect 68785 597 68831 643
rect 68909 597 68955 643
rect 69033 597 69079 643
rect 69157 597 69203 643
rect 69281 597 69327 643
rect 69405 597 69451 643
rect 69529 597 69575 643
rect 69653 597 69699 643
rect 69777 597 69823 643
rect 69901 597 69947 643
rect 70025 597 70071 643
rect 70149 597 70195 643
rect 70273 597 70319 643
rect 70397 597 70443 643
rect 70521 597 70567 643
rect 70645 597 70691 643
rect 70769 597 70815 643
rect 70893 597 70939 643
rect 71017 597 71063 643
rect 71141 597 71187 643
rect 71265 597 71311 643
rect 71389 597 71435 643
rect 71513 597 71559 643
rect 71637 597 71683 643
rect 71761 597 71807 643
rect 71885 597 71931 643
rect 72009 597 72055 643
rect 72133 597 72179 643
rect 72257 597 72303 643
rect 72381 597 72427 643
rect 72505 597 72551 643
rect 72629 597 72675 643
rect 72753 597 72799 643
rect 72877 597 72923 643
rect 73001 597 73047 643
rect 73125 597 73171 643
rect 73249 597 73295 643
rect 73373 597 73419 643
rect 73497 597 73543 643
rect 73621 597 73667 643
rect 73745 597 73791 643
rect 73869 597 73915 643
rect 73993 597 74039 643
rect 74117 597 74163 643
rect 74241 597 74287 643
rect 74365 597 74411 643
rect 74489 597 74535 643
rect 74613 597 74659 643
rect 74737 597 74783 643
rect 74861 597 74907 643
rect 74985 597 75031 643
rect 75109 597 75155 643
rect 75233 597 75279 643
rect 75357 597 75403 643
rect 75481 597 75527 643
rect 75605 597 75651 643
rect 75729 597 75775 643
rect 75853 597 75899 643
rect 75977 597 76023 643
rect 76101 597 76147 643
rect 76225 597 76271 643
rect 76349 597 76395 643
rect 76473 597 76519 643
rect 76597 597 76643 643
rect 76721 597 76767 643
rect 76845 597 76891 643
rect 76969 597 77015 643
rect 77093 597 77139 643
rect 77217 597 77263 643
rect 77341 597 77387 643
rect 77465 597 77511 643
rect 77589 597 77635 643
rect 77713 597 77759 643
rect 77837 597 77883 643
rect 77961 597 78007 643
rect 78085 597 78131 643
rect 78209 597 78255 643
rect 78333 597 78379 643
rect 78457 597 78503 643
rect 78581 597 78627 643
rect 78705 597 78751 643
rect 78829 597 78875 643
rect 78953 597 78999 643
rect 79077 597 79123 643
rect 79201 597 79247 643
rect 79325 597 79371 643
rect 79449 597 79495 643
rect 79573 597 79619 643
rect 79697 597 79743 643
rect 79821 597 79867 643
rect 79945 597 79991 643
rect 80069 597 80115 643
rect 80193 597 80239 643
rect 80317 597 80363 643
rect 80441 597 80487 643
rect 80565 597 80611 643
rect 80689 597 80735 643
rect 80813 597 80859 643
rect 80937 597 80983 643
rect 81061 597 81107 643
rect 81185 597 81231 643
rect 81309 597 81355 643
rect 81433 597 81479 643
rect 81557 597 81603 643
rect 81681 597 81727 643
rect 81805 597 81851 643
rect 81929 597 81975 643
rect 82053 597 82099 643
rect 82177 597 82223 643
rect 82301 597 82347 643
rect 82425 597 82471 643
rect 82549 597 82595 643
rect 82673 597 82719 643
rect 82797 597 82843 643
rect 82921 597 82967 643
rect 83045 597 83091 643
rect 83169 597 83215 643
rect 83293 597 83339 643
rect 83417 597 83463 643
rect 83541 597 83587 643
rect 83665 597 83711 643
rect 83789 597 83835 643
rect 83913 597 83959 643
rect 84037 597 84083 643
rect 84161 597 84207 643
rect 84285 597 84331 643
rect 84409 597 84455 643
rect 84533 597 84579 643
rect 84657 597 84703 643
rect 84781 597 84827 643
rect 84905 597 84951 643
rect 85029 597 85075 643
rect 85153 597 85199 643
rect 85277 597 85323 643
rect 85401 597 85447 643
rect 85525 597 85571 643
rect 85649 597 85695 643
<< metal1 >>
rect 0 67883 85808 67894
rect 0 67837 89 67883
rect 135 67837 213 67883
rect 259 67837 337 67883
rect 383 67837 461 67883
rect 507 67837 585 67883
rect 631 67837 709 67883
rect 755 67837 833 67883
rect 879 67837 957 67883
rect 1003 67837 1081 67883
rect 1127 67837 1205 67883
rect 1251 67837 1329 67883
rect 1375 67837 1453 67883
rect 1499 67837 1577 67883
rect 1623 67837 1701 67883
rect 1747 67837 1825 67883
rect 1871 67837 1949 67883
rect 1995 67837 2073 67883
rect 2119 67837 2197 67883
rect 2243 67837 2321 67883
rect 2367 67837 2445 67883
rect 2491 67837 2569 67883
rect 2615 67837 2693 67883
rect 2739 67837 2817 67883
rect 2863 67837 2941 67883
rect 2987 67837 3065 67883
rect 3111 67837 3189 67883
rect 3235 67837 3313 67883
rect 3359 67837 3437 67883
rect 3483 67837 3561 67883
rect 3607 67837 3685 67883
rect 3731 67837 3809 67883
rect 3855 67837 3933 67883
rect 3979 67837 4057 67883
rect 4103 67837 4181 67883
rect 4227 67837 4305 67883
rect 4351 67837 4429 67883
rect 4475 67837 4553 67883
rect 4599 67837 4677 67883
rect 4723 67837 4801 67883
rect 4847 67837 4925 67883
rect 4971 67837 5049 67883
rect 5095 67837 5173 67883
rect 5219 67837 5297 67883
rect 5343 67837 5421 67883
rect 5467 67837 5545 67883
rect 5591 67837 5669 67883
rect 5715 67837 5793 67883
rect 5839 67837 5917 67883
rect 5963 67837 6041 67883
rect 6087 67837 6165 67883
rect 6211 67837 6289 67883
rect 6335 67837 6413 67883
rect 6459 67837 6537 67883
rect 6583 67837 6661 67883
rect 6707 67837 6785 67883
rect 6831 67837 6909 67883
rect 6955 67837 7033 67883
rect 7079 67837 7157 67883
rect 7203 67837 7281 67883
rect 7327 67837 7405 67883
rect 7451 67837 7529 67883
rect 7575 67837 7653 67883
rect 7699 67837 7777 67883
rect 7823 67837 7901 67883
rect 7947 67837 8025 67883
rect 8071 67837 8149 67883
rect 8195 67837 8273 67883
rect 8319 67837 8397 67883
rect 8443 67837 8521 67883
rect 8567 67837 8645 67883
rect 8691 67837 8769 67883
rect 8815 67837 8893 67883
rect 8939 67837 9017 67883
rect 9063 67837 9141 67883
rect 9187 67837 9265 67883
rect 9311 67837 9389 67883
rect 9435 67837 9513 67883
rect 9559 67837 9637 67883
rect 9683 67837 9761 67883
rect 9807 67837 9885 67883
rect 9931 67837 10009 67883
rect 10055 67837 10133 67883
rect 10179 67837 10257 67883
rect 10303 67837 10381 67883
rect 10427 67837 10505 67883
rect 10551 67837 10629 67883
rect 10675 67837 10753 67883
rect 10799 67837 10877 67883
rect 10923 67837 11001 67883
rect 11047 67837 11125 67883
rect 11171 67837 11249 67883
rect 11295 67837 11373 67883
rect 11419 67837 11497 67883
rect 11543 67837 11621 67883
rect 11667 67837 11745 67883
rect 11791 67837 11869 67883
rect 11915 67837 11993 67883
rect 12039 67837 12117 67883
rect 12163 67837 12241 67883
rect 12287 67837 12365 67883
rect 12411 67837 12489 67883
rect 12535 67837 12613 67883
rect 12659 67837 12737 67883
rect 12783 67837 12861 67883
rect 12907 67837 12985 67883
rect 13031 67837 13109 67883
rect 13155 67837 13233 67883
rect 13279 67837 13357 67883
rect 13403 67837 13481 67883
rect 13527 67837 13605 67883
rect 13651 67837 13729 67883
rect 13775 67837 13853 67883
rect 13899 67837 13977 67883
rect 14023 67837 14101 67883
rect 14147 67837 14225 67883
rect 14271 67837 14349 67883
rect 14395 67837 14473 67883
rect 14519 67837 14597 67883
rect 14643 67837 14721 67883
rect 14767 67837 14845 67883
rect 14891 67837 14969 67883
rect 15015 67837 15093 67883
rect 15139 67837 15217 67883
rect 15263 67837 15341 67883
rect 15387 67837 15465 67883
rect 15511 67837 15589 67883
rect 15635 67837 15713 67883
rect 15759 67837 15837 67883
rect 15883 67837 15961 67883
rect 16007 67837 16085 67883
rect 16131 67837 16209 67883
rect 16255 67837 16333 67883
rect 16379 67837 16457 67883
rect 16503 67837 16581 67883
rect 16627 67837 16705 67883
rect 16751 67837 16829 67883
rect 16875 67837 16953 67883
rect 16999 67837 17077 67883
rect 17123 67837 17201 67883
rect 17247 67837 17325 67883
rect 17371 67837 17449 67883
rect 17495 67837 17573 67883
rect 17619 67837 17697 67883
rect 17743 67837 17821 67883
rect 17867 67837 17945 67883
rect 17991 67837 18069 67883
rect 18115 67837 18193 67883
rect 18239 67837 18317 67883
rect 18363 67837 18441 67883
rect 18487 67837 18565 67883
rect 18611 67837 18689 67883
rect 18735 67837 18813 67883
rect 18859 67837 18937 67883
rect 18983 67837 19061 67883
rect 19107 67837 19185 67883
rect 19231 67837 19309 67883
rect 19355 67837 19433 67883
rect 19479 67837 19557 67883
rect 19603 67837 19681 67883
rect 19727 67837 19805 67883
rect 19851 67837 19929 67883
rect 19975 67837 20053 67883
rect 20099 67837 20177 67883
rect 20223 67837 20301 67883
rect 20347 67837 20425 67883
rect 20471 67837 20549 67883
rect 20595 67837 20673 67883
rect 20719 67837 20797 67883
rect 20843 67837 20921 67883
rect 20967 67837 21045 67883
rect 21091 67837 21169 67883
rect 21215 67837 21293 67883
rect 21339 67837 21417 67883
rect 21463 67837 21541 67883
rect 21587 67837 21665 67883
rect 21711 67837 21789 67883
rect 21835 67837 21913 67883
rect 21959 67837 22037 67883
rect 22083 67837 22161 67883
rect 22207 67837 22285 67883
rect 22331 67837 22409 67883
rect 22455 67837 22533 67883
rect 22579 67837 22657 67883
rect 22703 67837 22781 67883
rect 22827 67837 22905 67883
rect 22951 67837 23029 67883
rect 23075 67837 23153 67883
rect 23199 67837 23277 67883
rect 23323 67837 23401 67883
rect 23447 67837 23525 67883
rect 23571 67837 23649 67883
rect 23695 67837 23773 67883
rect 23819 67837 23897 67883
rect 23943 67837 24021 67883
rect 24067 67837 24145 67883
rect 24191 67837 24269 67883
rect 24315 67837 24393 67883
rect 24439 67837 24517 67883
rect 24563 67837 24641 67883
rect 24687 67837 24765 67883
rect 24811 67837 24889 67883
rect 24935 67837 25013 67883
rect 25059 67837 25137 67883
rect 25183 67837 25261 67883
rect 25307 67837 25385 67883
rect 25431 67837 25509 67883
rect 25555 67837 25633 67883
rect 25679 67837 25757 67883
rect 25803 67837 25881 67883
rect 25927 67837 26005 67883
rect 26051 67837 26129 67883
rect 26175 67837 26253 67883
rect 26299 67837 26377 67883
rect 26423 67837 26501 67883
rect 26547 67837 26625 67883
rect 26671 67837 26749 67883
rect 26795 67837 26873 67883
rect 26919 67837 26997 67883
rect 27043 67837 27121 67883
rect 27167 67837 27245 67883
rect 27291 67837 27369 67883
rect 27415 67837 27493 67883
rect 27539 67837 27617 67883
rect 27663 67837 27741 67883
rect 27787 67837 27865 67883
rect 27911 67837 27989 67883
rect 28035 67837 28113 67883
rect 28159 67837 28237 67883
rect 28283 67837 28361 67883
rect 28407 67837 28485 67883
rect 28531 67837 28609 67883
rect 28655 67837 28733 67883
rect 28779 67837 28857 67883
rect 28903 67837 28981 67883
rect 29027 67837 29105 67883
rect 29151 67837 29229 67883
rect 29275 67837 29353 67883
rect 29399 67837 29477 67883
rect 29523 67837 29601 67883
rect 29647 67837 29725 67883
rect 29771 67837 29849 67883
rect 29895 67837 29973 67883
rect 30019 67837 30097 67883
rect 30143 67837 30221 67883
rect 30267 67837 30345 67883
rect 30391 67837 30469 67883
rect 30515 67837 30593 67883
rect 30639 67837 30717 67883
rect 30763 67837 30841 67883
rect 30887 67837 30965 67883
rect 31011 67837 31089 67883
rect 31135 67837 31213 67883
rect 31259 67837 31337 67883
rect 31383 67837 31461 67883
rect 31507 67837 31585 67883
rect 31631 67837 31709 67883
rect 31755 67837 31833 67883
rect 31879 67837 31957 67883
rect 32003 67837 32081 67883
rect 32127 67837 32205 67883
rect 32251 67837 32329 67883
rect 32375 67837 32453 67883
rect 32499 67837 32577 67883
rect 32623 67837 32701 67883
rect 32747 67837 32825 67883
rect 32871 67837 32949 67883
rect 32995 67837 33073 67883
rect 33119 67837 33197 67883
rect 33243 67837 33321 67883
rect 33367 67837 33445 67883
rect 33491 67837 33569 67883
rect 33615 67837 33693 67883
rect 33739 67837 33817 67883
rect 33863 67837 33941 67883
rect 33987 67837 34065 67883
rect 34111 67837 34189 67883
rect 34235 67837 34313 67883
rect 34359 67837 34437 67883
rect 34483 67837 34561 67883
rect 34607 67837 34685 67883
rect 34731 67837 34809 67883
rect 34855 67837 34933 67883
rect 34979 67837 35057 67883
rect 35103 67837 35181 67883
rect 35227 67837 35305 67883
rect 35351 67837 35429 67883
rect 35475 67837 35553 67883
rect 35599 67837 35677 67883
rect 35723 67837 35801 67883
rect 35847 67837 35925 67883
rect 35971 67837 36049 67883
rect 36095 67837 36173 67883
rect 36219 67837 36297 67883
rect 36343 67837 36421 67883
rect 36467 67837 36545 67883
rect 36591 67837 36669 67883
rect 36715 67837 36793 67883
rect 36839 67837 36917 67883
rect 36963 67837 37041 67883
rect 37087 67837 37165 67883
rect 37211 67837 37289 67883
rect 37335 67837 37413 67883
rect 37459 67837 37537 67883
rect 37583 67837 37661 67883
rect 37707 67837 37785 67883
rect 37831 67837 37909 67883
rect 37955 67837 38033 67883
rect 38079 67837 38157 67883
rect 38203 67837 38281 67883
rect 38327 67837 38405 67883
rect 38451 67837 38529 67883
rect 38575 67837 38653 67883
rect 38699 67837 38777 67883
rect 38823 67837 38901 67883
rect 38947 67837 39025 67883
rect 39071 67837 39149 67883
rect 39195 67837 39273 67883
rect 39319 67837 39397 67883
rect 39443 67837 39521 67883
rect 39567 67837 39645 67883
rect 39691 67837 39769 67883
rect 39815 67837 39893 67883
rect 39939 67837 40017 67883
rect 40063 67837 40141 67883
rect 40187 67837 40265 67883
rect 40311 67837 40389 67883
rect 40435 67837 40513 67883
rect 40559 67837 40637 67883
rect 40683 67837 40761 67883
rect 40807 67837 40885 67883
rect 40931 67837 41009 67883
rect 41055 67837 41133 67883
rect 41179 67837 41257 67883
rect 41303 67837 41381 67883
rect 41427 67837 41505 67883
rect 41551 67837 41629 67883
rect 41675 67837 41753 67883
rect 41799 67837 41877 67883
rect 41923 67837 42001 67883
rect 42047 67837 42125 67883
rect 42171 67837 42249 67883
rect 42295 67837 42373 67883
rect 42419 67837 42497 67883
rect 42543 67837 42621 67883
rect 42667 67837 42745 67883
rect 42791 67837 42869 67883
rect 42915 67837 42993 67883
rect 43039 67837 43117 67883
rect 43163 67837 43241 67883
rect 43287 67837 43365 67883
rect 43411 67837 43489 67883
rect 43535 67837 43613 67883
rect 43659 67837 43737 67883
rect 43783 67837 43861 67883
rect 43907 67837 43985 67883
rect 44031 67837 44109 67883
rect 44155 67837 44233 67883
rect 44279 67837 44357 67883
rect 44403 67837 44481 67883
rect 44527 67837 44605 67883
rect 44651 67837 44729 67883
rect 44775 67837 44853 67883
rect 44899 67837 44977 67883
rect 45023 67837 45101 67883
rect 45147 67837 45225 67883
rect 45271 67837 45349 67883
rect 45395 67837 45473 67883
rect 45519 67837 45597 67883
rect 45643 67837 45721 67883
rect 45767 67837 45845 67883
rect 45891 67837 45969 67883
rect 46015 67837 46093 67883
rect 46139 67837 46217 67883
rect 46263 67837 46341 67883
rect 46387 67837 46465 67883
rect 46511 67837 46589 67883
rect 46635 67837 46713 67883
rect 46759 67837 46837 67883
rect 46883 67837 46961 67883
rect 47007 67837 47085 67883
rect 47131 67837 47209 67883
rect 47255 67837 47333 67883
rect 47379 67837 47457 67883
rect 47503 67837 47581 67883
rect 47627 67837 47705 67883
rect 47751 67837 47829 67883
rect 47875 67837 47953 67883
rect 47999 67837 48077 67883
rect 48123 67837 48201 67883
rect 48247 67837 48325 67883
rect 48371 67837 48449 67883
rect 48495 67837 48573 67883
rect 48619 67837 48697 67883
rect 48743 67837 48821 67883
rect 48867 67837 48945 67883
rect 48991 67837 49069 67883
rect 49115 67837 49193 67883
rect 49239 67837 49317 67883
rect 49363 67837 49441 67883
rect 49487 67837 49565 67883
rect 49611 67837 49689 67883
rect 49735 67837 49813 67883
rect 49859 67837 49937 67883
rect 49983 67837 50061 67883
rect 50107 67837 50185 67883
rect 50231 67837 50309 67883
rect 50355 67837 50433 67883
rect 50479 67837 50557 67883
rect 50603 67837 50681 67883
rect 50727 67837 50805 67883
rect 50851 67837 50929 67883
rect 50975 67837 51053 67883
rect 51099 67837 51177 67883
rect 51223 67837 51301 67883
rect 51347 67837 51425 67883
rect 51471 67837 51549 67883
rect 51595 67837 51673 67883
rect 51719 67837 51797 67883
rect 51843 67837 51921 67883
rect 51967 67837 52045 67883
rect 52091 67837 52169 67883
rect 52215 67837 52293 67883
rect 52339 67837 52417 67883
rect 52463 67837 52541 67883
rect 52587 67837 52665 67883
rect 52711 67837 52789 67883
rect 52835 67837 52913 67883
rect 52959 67837 53037 67883
rect 53083 67837 53161 67883
rect 53207 67837 53285 67883
rect 53331 67837 53409 67883
rect 53455 67837 53533 67883
rect 53579 67837 53657 67883
rect 53703 67837 53781 67883
rect 53827 67837 53905 67883
rect 53951 67837 54029 67883
rect 54075 67837 54153 67883
rect 54199 67837 54277 67883
rect 54323 67837 54401 67883
rect 54447 67837 54525 67883
rect 54571 67837 54649 67883
rect 54695 67837 54773 67883
rect 54819 67837 54897 67883
rect 54943 67837 55021 67883
rect 55067 67837 55145 67883
rect 55191 67837 55269 67883
rect 55315 67837 55393 67883
rect 55439 67837 55517 67883
rect 55563 67837 55641 67883
rect 55687 67837 55765 67883
rect 55811 67837 55889 67883
rect 55935 67837 56013 67883
rect 56059 67837 56137 67883
rect 56183 67837 56261 67883
rect 56307 67837 56385 67883
rect 56431 67837 56509 67883
rect 56555 67837 56633 67883
rect 56679 67837 56757 67883
rect 56803 67837 56881 67883
rect 56927 67837 57005 67883
rect 57051 67837 57129 67883
rect 57175 67837 57253 67883
rect 57299 67837 57377 67883
rect 57423 67837 57501 67883
rect 57547 67837 57625 67883
rect 57671 67837 57749 67883
rect 57795 67837 57873 67883
rect 57919 67837 57997 67883
rect 58043 67837 58121 67883
rect 58167 67837 58245 67883
rect 58291 67837 58369 67883
rect 58415 67837 58493 67883
rect 58539 67837 58617 67883
rect 58663 67837 58741 67883
rect 58787 67837 58865 67883
rect 58911 67837 58989 67883
rect 59035 67837 59113 67883
rect 59159 67837 59237 67883
rect 59283 67837 59361 67883
rect 59407 67837 59485 67883
rect 59531 67837 59609 67883
rect 59655 67837 59733 67883
rect 59779 67837 59857 67883
rect 59903 67837 59981 67883
rect 60027 67837 60105 67883
rect 60151 67837 60229 67883
rect 60275 67837 60353 67883
rect 60399 67837 60477 67883
rect 60523 67837 60601 67883
rect 60647 67837 60725 67883
rect 60771 67837 60849 67883
rect 60895 67837 60973 67883
rect 61019 67837 61097 67883
rect 61143 67837 61221 67883
rect 61267 67837 61345 67883
rect 61391 67837 61469 67883
rect 61515 67837 61593 67883
rect 61639 67837 61717 67883
rect 61763 67837 61841 67883
rect 61887 67837 61965 67883
rect 62011 67837 62089 67883
rect 62135 67837 62213 67883
rect 62259 67837 62337 67883
rect 62383 67837 62461 67883
rect 62507 67837 62585 67883
rect 62631 67837 62709 67883
rect 62755 67837 62833 67883
rect 62879 67837 62957 67883
rect 63003 67837 63081 67883
rect 63127 67837 63205 67883
rect 63251 67837 63329 67883
rect 63375 67837 63453 67883
rect 63499 67837 63577 67883
rect 63623 67837 63701 67883
rect 63747 67837 63825 67883
rect 63871 67837 63949 67883
rect 63995 67837 64073 67883
rect 64119 67837 64197 67883
rect 64243 67837 64321 67883
rect 64367 67837 64445 67883
rect 64491 67837 64569 67883
rect 64615 67837 64693 67883
rect 64739 67837 64817 67883
rect 64863 67837 64941 67883
rect 64987 67837 65065 67883
rect 65111 67837 65189 67883
rect 65235 67837 65313 67883
rect 65359 67837 65437 67883
rect 65483 67837 65561 67883
rect 65607 67837 65685 67883
rect 65731 67837 65809 67883
rect 65855 67837 65933 67883
rect 65979 67837 66057 67883
rect 66103 67837 66181 67883
rect 66227 67837 66305 67883
rect 66351 67837 66429 67883
rect 66475 67837 66553 67883
rect 66599 67837 66677 67883
rect 66723 67837 66801 67883
rect 66847 67837 66925 67883
rect 66971 67837 67049 67883
rect 67095 67837 67173 67883
rect 67219 67837 67297 67883
rect 67343 67837 67421 67883
rect 67467 67837 67545 67883
rect 67591 67837 67669 67883
rect 67715 67837 67793 67883
rect 67839 67837 67917 67883
rect 67963 67837 68041 67883
rect 68087 67837 68165 67883
rect 68211 67837 68289 67883
rect 68335 67837 68413 67883
rect 68459 67837 68537 67883
rect 68583 67837 68661 67883
rect 68707 67837 68785 67883
rect 68831 67837 68909 67883
rect 68955 67837 69033 67883
rect 69079 67837 69157 67883
rect 69203 67837 69281 67883
rect 69327 67837 69405 67883
rect 69451 67837 69529 67883
rect 69575 67837 69653 67883
rect 69699 67837 69777 67883
rect 69823 67837 69901 67883
rect 69947 67837 70025 67883
rect 70071 67837 70149 67883
rect 70195 67837 70273 67883
rect 70319 67837 70397 67883
rect 70443 67837 70521 67883
rect 70567 67837 70645 67883
rect 70691 67837 70769 67883
rect 70815 67837 70893 67883
rect 70939 67837 71017 67883
rect 71063 67837 71141 67883
rect 71187 67837 71265 67883
rect 71311 67837 71389 67883
rect 71435 67837 71513 67883
rect 71559 67837 71637 67883
rect 71683 67837 71761 67883
rect 71807 67837 71885 67883
rect 71931 67837 72009 67883
rect 72055 67837 72133 67883
rect 72179 67837 72257 67883
rect 72303 67837 72381 67883
rect 72427 67837 72505 67883
rect 72551 67837 72629 67883
rect 72675 67837 72753 67883
rect 72799 67837 72877 67883
rect 72923 67837 73001 67883
rect 73047 67837 73125 67883
rect 73171 67837 73249 67883
rect 73295 67837 73373 67883
rect 73419 67837 73497 67883
rect 73543 67837 73621 67883
rect 73667 67837 73745 67883
rect 73791 67837 73869 67883
rect 73915 67837 73993 67883
rect 74039 67837 74117 67883
rect 74163 67837 74241 67883
rect 74287 67837 74365 67883
rect 74411 67837 74489 67883
rect 74535 67837 74613 67883
rect 74659 67837 74737 67883
rect 74783 67837 74861 67883
rect 74907 67837 74985 67883
rect 75031 67837 75109 67883
rect 75155 67837 75233 67883
rect 75279 67837 75357 67883
rect 75403 67837 75481 67883
rect 75527 67837 75605 67883
rect 75651 67837 75729 67883
rect 75775 67837 75853 67883
rect 75899 67837 75977 67883
rect 76023 67837 76101 67883
rect 76147 67837 76225 67883
rect 76271 67837 76349 67883
rect 76395 67837 76473 67883
rect 76519 67837 76597 67883
rect 76643 67837 76721 67883
rect 76767 67837 76845 67883
rect 76891 67837 76969 67883
rect 77015 67837 77093 67883
rect 77139 67837 77217 67883
rect 77263 67837 77341 67883
rect 77387 67837 77465 67883
rect 77511 67837 77589 67883
rect 77635 67837 77713 67883
rect 77759 67837 77837 67883
rect 77883 67837 77961 67883
rect 78007 67837 78085 67883
rect 78131 67837 78209 67883
rect 78255 67837 78333 67883
rect 78379 67837 78457 67883
rect 78503 67837 78581 67883
rect 78627 67837 78705 67883
rect 78751 67837 78829 67883
rect 78875 67837 78953 67883
rect 78999 67837 79077 67883
rect 79123 67837 79201 67883
rect 79247 67837 79325 67883
rect 79371 67837 79449 67883
rect 79495 67837 79573 67883
rect 79619 67837 79697 67883
rect 79743 67837 79821 67883
rect 79867 67837 79945 67883
rect 79991 67837 80069 67883
rect 80115 67837 80193 67883
rect 80239 67837 80317 67883
rect 80363 67837 80441 67883
rect 80487 67837 80565 67883
rect 80611 67837 80689 67883
rect 80735 67837 80813 67883
rect 80859 67837 80937 67883
rect 80983 67837 81061 67883
rect 81107 67837 81185 67883
rect 81231 67837 81309 67883
rect 81355 67837 81433 67883
rect 81479 67837 81557 67883
rect 81603 67837 81681 67883
rect 81727 67837 81805 67883
rect 81851 67837 81929 67883
rect 81975 67837 82053 67883
rect 82099 67837 82177 67883
rect 82223 67837 82301 67883
rect 82347 67837 82425 67883
rect 82471 67837 82549 67883
rect 82595 67837 82673 67883
rect 82719 67837 82797 67883
rect 82843 67837 82921 67883
rect 82967 67837 83045 67883
rect 83091 67837 83169 67883
rect 83215 67837 83293 67883
rect 83339 67837 83417 67883
rect 83463 67837 83541 67883
rect 83587 67837 83665 67883
rect 83711 67837 83789 67883
rect 83835 67837 83913 67883
rect 83959 67837 84037 67883
rect 84083 67837 84161 67883
rect 84207 67837 84285 67883
rect 84331 67837 84409 67883
rect 84455 67837 84533 67883
rect 84579 67837 84657 67883
rect 84703 67837 84781 67883
rect 84827 67837 84905 67883
rect 84951 67837 85029 67883
rect 85075 67837 85153 67883
rect 85199 67837 85277 67883
rect 85323 67837 85401 67883
rect 85447 67837 85525 67883
rect 85571 67837 85649 67883
rect 85695 67837 85808 67883
rect 0 67759 85808 67837
rect 0 67713 89 67759
rect 135 67713 213 67759
rect 259 67713 337 67759
rect 383 67713 461 67759
rect 507 67713 585 67759
rect 631 67713 709 67759
rect 755 67713 833 67759
rect 879 67713 957 67759
rect 1003 67713 1081 67759
rect 1127 67713 1205 67759
rect 1251 67713 1329 67759
rect 1375 67713 1453 67759
rect 1499 67713 1577 67759
rect 1623 67713 1701 67759
rect 1747 67713 1825 67759
rect 1871 67713 1949 67759
rect 1995 67713 2073 67759
rect 2119 67713 2197 67759
rect 2243 67713 2321 67759
rect 2367 67713 2445 67759
rect 2491 67713 2569 67759
rect 2615 67713 2693 67759
rect 2739 67713 2817 67759
rect 2863 67713 2941 67759
rect 2987 67713 3065 67759
rect 3111 67713 3189 67759
rect 3235 67713 3313 67759
rect 3359 67713 3437 67759
rect 3483 67713 3561 67759
rect 3607 67713 3685 67759
rect 3731 67713 3809 67759
rect 3855 67713 3933 67759
rect 3979 67713 4057 67759
rect 4103 67713 4181 67759
rect 4227 67713 4305 67759
rect 4351 67713 4429 67759
rect 4475 67713 4553 67759
rect 4599 67713 4677 67759
rect 4723 67713 4801 67759
rect 4847 67713 4925 67759
rect 4971 67713 5049 67759
rect 5095 67713 5173 67759
rect 5219 67713 5297 67759
rect 5343 67713 5421 67759
rect 5467 67713 5545 67759
rect 5591 67713 5669 67759
rect 5715 67713 5793 67759
rect 5839 67713 5917 67759
rect 5963 67713 6041 67759
rect 6087 67713 6165 67759
rect 6211 67713 6289 67759
rect 6335 67713 6413 67759
rect 6459 67713 6537 67759
rect 6583 67713 6661 67759
rect 6707 67713 6785 67759
rect 6831 67713 6909 67759
rect 6955 67713 7033 67759
rect 7079 67713 7157 67759
rect 7203 67713 7281 67759
rect 7327 67713 7405 67759
rect 7451 67713 7529 67759
rect 7575 67713 7653 67759
rect 7699 67713 7777 67759
rect 7823 67713 7901 67759
rect 7947 67713 8025 67759
rect 8071 67713 8149 67759
rect 8195 67713 8273 67759
rect 8319 67713 8397 67759
rect 8443 67713 8521 67759
rect 8567 67713 8645 67759
rect 8691 67713 8769 67759
rect 8815 67713 8893 67759
rect 8939 67713 9017 67759
rect 9063 67713 9141 67759
rect 9187 67713 9265 67759
rect 9311 67713 9389 67759
rect 9435 67713 9513 67759
rect 9559 67713 9637 67759
rect 9683 67713 9761 67759
rect 9807 67713 9885 67759
rect 9931 67713 10009 67759
rect 10055 67713 10133 67759
rect 10179 67713 10257 67759
rect 10303 67713 10381 67759
rect 10427 67713 10505 67759
rect 10551 67713 10629 67759
rect 10675 67713 10753 67759
rect 10799 67713 10877 67759
rect 10923 67713 11001 67759
rect 11047 67713 11125 67759
rect 11171 67713 11249 67759
rect 11295 67713 11373 67759
rect 11419 67713 11497 67759
rect 11543 67713 11621 67759
rect 11667 67713 11745 67759
rect 11791 67713 11869 67759
rect 11915 67713 11993 67759
rect 12039 67713 12117 67759
rect 12163 67713 12241 67759
rect 12287 67713 12365 67759
rect 12411 67713 12489 67759
rect 12535 67713 12613 67759
rect 12659 67713 12737 67759
rect 12783 67713 12861 67759
rect 12907 67713 12985 67759
rect 13031 67713 13109 67759
rect 13155 67713 13233 67759
rect 13279 67713 13357 67759
rect 13403 67713 13481 67759
rect 13527 67713 13605 67759
rect 13651 67713 13729 67759
rect 13775 67713 13853 67759
rect 13899 67713 13977 67759
rect 14023 67713 14101 67759
rect 14147 67713 14225 67759
rect 14271 67713 14349 67759
rect 14395 67713 14473 67759
rect 14519 67713 14597 67759
rect 14643 67713 14721 67759
rect 14767 67713 14845 67759
rect 14891 67713 14969 67759
rect 15015 67713 15093 67759
rect 15139 67713 15217 67759
rect 15263 67713 15341 67759
rect 15387 67713 15465 67759
rect 15511 67713 15589 67759
rect 15635 67713 15713 67759
rect 15759 67713 15837 67759
rect 15883 67713 15961 67759
rect 16007 67713 16085 67759
rect 16131 67713 16209 67759
rect 16255 67713 16333 67759
rect 16379 67713 16457 67759
rect 16503 67713 16581 67759
rect 16627 67713 16705 67759
rect 16751 67713 16829 67759
rect 16875 67713 16953 67759
rect 16999 67713 17077 67759
rect 17123 67713 17201 67759
rect 17247 67713 17325 67759
rect 17371 67713 17449 67759
rect 17495 67713 17573 67759
rect 17619 67713 17697 67759
rect 17743 67713 17821 67759
rect 17867 67713 17945 67759
rect 17991 67713 18069 67759
rect 18115 67713 18193 67759
rect 18239 67713 18317 67759
rect 18363 67713 18441 67759
rect 18487 67713 18565 67759
rect 18611 67713 18689 67759
rect 18735 67713 18813 67759
rect 18859 67713 18937 67759
rect 18983 67713 19061 67759
rect 19107 67713 19185 67759
rect 19231 67713 19309 67759
rect 19355 67713 19433 67759
rect 19479 67713 19557 67759
rect 19603 67713 19681 67759
rect 19727 67713 19805 67759
rect 19851 67713 19929 67759
rect 19975 67713 20053 67759
rect 20099 67713 20177 67759
rect 20223 67713 20301 67759
rect 20347 67713 20425 67759
rect 20471 67713 20549 67759
rect 20595 67713 20673 67759
rect 20719 67713 20797 67759
rect 20843 67713 20921 67759
rect 20967 67713 21045 67759
rect 21091 67713 21169 67759
rect 21215 67713 21293 67759
rect 21339 67713 21417 67759
rect 21463 67713 21541 67759
rect 21587 67713 21665 67759
rect 21711 67713 21789 67759
rect 21835 67713 21913 67759
rect 21959 67713 22037 67759
rect 22083 67713 22161 67759
rect 22207 67713 22285 67759
rect 22331 67713 22409 67759
rect 22455 67713 22533 67759
rect 22579 67713 22657 67759
rect 22703 67713 22781 67759
rect 22827 67713 22905 67759
rect 22951 67713 23029 67759
rect 23075 67713 23153 67759
rect 23199 67713 23277 67759
rect 23323 67713 23401 67759
rect 23447 67713 23525 67759
rect 23571 67713 23649 67759
rect 23695 67713 23773 67759
rect 23819 67713 23897 67759
rect 23943 67713 24021 67759
rect 24067 67713 24145 67759
rect 24191 67713 24269 67759
rect 24315 67713 24393 67759
rect 24439 67713 24517 67759
rect 24563 67713 24641 67759
rect 24687 67713 24765 67759
rect 24811 67713 24889 67759
rect 24935 67713 25013 67759
rect 25059 67713 25137 67759
rect 25183 67713 25261 67759
rect 25307 67713 25385 67759
rect 25431 67713 25509 67759
rect 25555 67713 25633 67759
rect 25679 67713 25757 67759
rect 25803 67713 25881 67759
rect 25927 67713 26005 67759
rect 26051 67713 26129 67759
rect 26175 67713 26253 67759
rect 26299 67713 26377 67759
rect 26423 67713 26501 67759
rect 26547 67713 26625 67759
rect 26671 67713 26749 67759
rect 26795 67713 26873 67759
rect 26919 67713 26997 67759
rect 27043 67713 27121 67759
rect 27167 67713 27245 67759
rect 27291 67713 27369 67759
rect 27415 67713 27493 67759
rect 27539 67713 27617 67759
rect 27663 67713 27741 67759
rect 27787 67713 27865 67759
rect 27911 67713 27989 67759
rect 28035 67713 28113 67759
rect 28159 67713 28237 67759
rect 28283 67713 28361 67759
rect 28407 67713 28485 67759
rect 28531 67713 28609 67759
rect 28655 67713 28733 67759
rect 28779 67713 28857 67759
rect 28903 67713 28981 67759
rect 29027 67713 29105 67759
rect 29151 67713 29229 67759
rect 29275 67713 29353 67759
rect 29399 67713 29477 67759
rect 29523 67713 29601 67759
rect 29647 67713 29725 67759
rect 29771 67713 29849 67759
rect 29895 67713 29973 67759
rect 30019 67713 30097 67759
rect 30143 67713 30221 67759
rect 30267 67713 30345 67759
rect 30391 67713 30469 67759
rect 30515 67713 30593 67759
rect 30639 67713 30717 67759
rect 30763 67713 30841 67759
rect 30887 67713 30965 67759
rect 31011 67713 31089 67759
rect 31135 67713 31213 67759
rect 31259 67713 31337 67759
rect 31383 67713 31461 67759
rect 31507 67713 31585 67759
rect 31631 67713 31709 67759
rect 31755 67713 31833 67759
rect 31879 67713 31957 67759
rect 32003 67713 32081 67759
rect 32127 67713 32205 67759
rect 32251 67713 32329 67759
rect 32375 67713 32453 67759
rect 32499 67713 32577 67759
rect 32623 67713 32701 67759
rect 32747 67713 32825 67759
rect 32871 67713 32949 67759
rect 32995 67713 33073 67759
rect 33119 67713 33197 67759
rect 33243 67713 33321 67759
rect 33367 67713 33445 67759
rect 33491 67713 33569 67759
rect 33615 67713 33693 67759
rect 33739 67713 33817 67759
rect 33863 67713 33941 67759
rect 33987 67713 34065 67759
rect 34111 67713 34189 67759
rect 34235 67713 34313 67759
rect 34359 67713 34437 67759
rect 34483 67713 34561 67759
rect 34607 67713 34685 67759
rect 34731 67713 34809 67759
rect 34855 67713 34933 67759
rect 34979 67713 35057 67759
rect 35103 67713 35181 67759
rect 35227 67713 35305 67759
rect 35351 67713 35429 67759
rect 35475 67713 35553 67759
rect 35599 67713 35677 67759
rect 35723 67713 35801 67759
rect 35847 67713 35925 67759
rect 35971 67713 36049 67759
rect 36095 67713 36173 67759
rect 36219 67713 36297 67759
rect 36343 67713 36421 67759
rect 36467 67713 36545 67759
rect 36591 67713 36669 67759
rect 36715 67713 36793 67759
rect 36839 67713 36917 67759
rect 36963 67713 37041 67759
rect 37087 67713 37165 67759
rect 37211 67713 37289 67759
rect 37335 67713 37413 67759
rect 37459 67713 37537 67759
rect 37583 67713 37661 67759
rect 37707 67713 37785 67759
rect 37831 67713 37909 67759
rect 37955 67713 38033 67759
rect 38079 67713 38157 67759
rect 38203 67713 38281 67759
rect 38327 67713 38405 67759
rect 38451 67713 38529 67759
rect 38575 67713 38653 67759
rect 38699 67713 38777 67759
rect 38823 67713 38901 67759
rect 38947 67713 39025 67759
rect 39071 67713 39149 67759
rect 39195 67713 39273 67759
rect 39319 67713 39397 67759
rect 39443 67713 39521 67759
rect 39567 67713 39645 67759
rect 39691 67713 39769 67759
rect 39815 67713 39893 67759
rect 39939 67713 40017 67759
rect 40063 67713 40141 67759
rect 40187 67713 40265 67759
rect 40311 67713 40389 67759
rect 40435 67713 40513 67759
rect 40559 67713 40637 67759
rect 40683 67713 40761 67759
rect 40807 67713 40885 67759
rect 40931 67713 41009 67759
rect 41055 67713 41133 67759
rect 41179 67713 41257 67759
rect 41303 67713 41381 67759
rect 41427 67713 41505 67759
rect 41551 67713 41629 67759
rect 41675 67713 41753 67759
rect 41799 67713 41877 67759
rect 41923 67713 42001 67759
rect 42047 67713 42125 67759
rect 42171 67713 42249 67759
rect 42295 67713 42373 67759
rect 42419 67713 42497 67759
rect 42543 67713 42621 67759
rect 42667 67713 42745 67759
rect 42791 67713 42869 67759
rect 42915 67713 42993 67759
rect 43039 67713 43117 67759
rect 43163 67713 43241 67759
rect 43287 67713 43365 67759
rect 43411 67713 43489 67759
rect 43535 67713 43613 67759
rect 43659 67713 43737 67759
rect 43783 67713 43861 67759
rect 43907 67713 43985 67759
rect 44031 67713 44109 67759
rect 44155 67713 44233 67759
rect 44279 67713 44357 67759
rect 44403 67713 44481 67759
rect 44527 67713 44605 67759
rect 44651 67713 44729 67759
rect 44775 67713 44853 67759
rect 44899 67713 44977 67759
rect 45023 67713 45101 67759
rect 45147 67713 45225 67759
rect 45271 67713 45349 67759
rect 45395 67713 45473 67759
rect 45519 67713 45597 67759
rect 45643 67713 45721 67759
rect 45767 67713 45845 67759
rect 45891 67713 45969 67759
rect 46015 67713 46093 67759
rect 46139 67713 46217 67759
rect 46263 67713 46341 67759
rect 46387 67713 46465 67759
rect 46511 67713 46589 67759
rect 46635 67713 46713 67759
rect 46759 67713 46837 67759
rect 46883 67713 46961 67759
rect 47007 67713 47085 67759
rect 47131 67713 47209 67759
rect 47255 67713 47333 67759
rect 47379 67713 47457 67759
rect 47503 67713 47581 67759
rect 47627 67713 47705 67759
rect 47751 67713 47829 67759
rect 47875 67713 47953 67759
rect 47999 67713 48077 67759
rect 48123 67713 48201 67759
rect 48247 67713 48325 67759
rect 48371 67713 48449 67759
rect 48495 67713 48573 67759
rect 48619 67713 48697 67759
rect 48743 67713 48821 67759
rect 48867 67713 48945 67759
rect 48991 67713 49069 67759
rect 49115 67713 49193 67759
rect 49239 67713 49317 67759
rect 49363 67713 49441 67759
rect 49487 67713 49565 67759
rect 49611 67713 49689 67759
rect 49735 67713 49813 67759
rect 49859 67713 49937 67759
rect 49983 67713 50061 67759
rect 50107 67713 50185 67759
rect 50231 67713 50309 67759
rect 50355 67713 50433 67759
rect 50479 67713 50557 67759
rect 50603 67713 50681 67759
rect 50727 67713 50805 67759
rect 50851 67713 50929 67759
rect 50975 67713 51053 67759
rect 51099 67713 51177 67759
rect 51223 67713 51301 67759
rect 51347 67713 51425 67759
rect 51471 67713 51549 67759
rect 51595 67713 51673 67759
rect 51719 67713 51797 67759
rect 51843 67713 51921 67759
rect 51967 67713 52045 67759
rect 52091 67713 52169 67759
rect 52215 67713 52293 67759
rect 52339 67713 52417 67759
rect 52463 67713 52541 67759
rect 52587 67713 52665 67759
rect 52711 67713 52789 67759
rect 52835 67713 52913 67759
rect 52959 67713 53037 67759
rect 53083 67713 53161 67759
rect 53207 67713 53285 67759
rect 53331 67713 53409 67759
rect 53455 67713 53533 67759
rect 53579 67713 53657 67759
rect 53703 67713 53781 67759
rect 53827 67713 53905 67759
rect 53951 67713 54029 67759
rect 54075 67713 54153 67759
rect 54199 67713 54277 67759
rect 54323 67713 54401 67759
rect 54447 67713 54525 67759
rect 54571 67713 54649 67759
rect 54695 67713 54773 67759
rect 54819 67713 54897 67759
rect 54943 67713 55021 67759
rect 55067 67713 55145 67759
rect 55191 67713 55269 67759
rect 55315 67713 55393 67759
rect 55439 67713 55517 67759
rect 55563 67713 55641 67759
rect 55687 67713 55765 67759
rect 55811 67713 55889 67759
rect 55935 67713 56013 67759
rect 56059 67713 56137 67759
rect 56183 67713 56261 67759
rect 56307 67713 56385 67759
rect 56431 67713 56509 67759
rect 56555 67713 56633 67759
rect 56679 67713 56757 67759
rect 56803 67713 56881 67759
rect 56927 67713 57005 67759
rect 57051 67713 57129 67759
rect 57175 67713 57253 67759
rect 57299 67713 57377 67759
rect 57423 67713 57501 67759
rect 57547 67713 57625 67759
rect 57671 67713 57749 67759
rect 57795 67713 57873 67759
rect 57919 67713 57997 67759
rect 58043 67713 58121 67759
rect 58167 67713 58245 67759
rect 58291 67713 58369 67759
rect 58415 67713 58493 67759
rect 58539 67713 58617 67759
rect 58663 67713 58741 67759
rect 58787 67713 58865 67759
rect 58911 67713 58989 67759
rect 59035 67713 59113 67759
rect 59159 67713 59237 67759
rect 59283 67713 59361 67759
rect 59407 67713 59485 67759
rect 59531 67713 59609 67759
rect 59655 67713 59733 67759
rect 59779 67713 59857 67759
rect 59903 67713 59981 67759
rect 60027 67713 60105 67759
rect 60151 67713 60229 67759
rect 60275 67713 60353 67759
rect 60399 67713 60477 67759
rect 60523 67713 60601 67759
rect 60647 67713 60725 67759
rect 60771 67713 60849 67759
rect 60895 67713 60973 67759
rect 61019 67713 61097 67759
rect 61143 67713 61221 67759
rect 61267 67713 61345 67759
rect 61391 67713 61469 67759
rect 61515 67713 61593 67759
rect 61639 67713 61717 67759
rect 61763 67713 61841 67759
rect 61887 67713 61965 67759
rect 62011 67713 62089 67759
rect 62135 67713 62213 67759
rect 62259 67713 62337 67759
rect 62383 67713 62461 67759
rect 62507 67713 62585 67759
rect 62631 67713 62709 67759
rect 62755 67713 62833 67759
rect 62879 67713 62957 67759
rect 63003 67713 63081 67759
rect 63127 67713 63205 67759
rect 63251 67713 63329 67759
rect 63375 67713 63453 67759
rect 63499 67713 63577 67759
rect 63623 67713 63701 67759
rect 63747 67713 63825 67759
rect 63871 67713 63949 67759
rect 63995 67713 64073 67759
rect 64119 67713 64197 67759
rect 64243 67713 64321 67759
rect 64367 67713 64445 67759
rect 64491 67713 64569 67759
rect 64615 67713 64693 67759
rect 64739 67713 64817 67759
rect 64863 67713 64941 67759
rect 64987 67713 65065 67759
rect 65111 67713 65189 67759
rect 65235 67713 65313 67759
rect 65359 67713 65437 67759
rect 65483 67713 65561 67759
rect 65607 67713 65685 67759
rect 65731 67713 65809 67759
rect 65855 67713 65933 67759
rect 65979 67713 66057 67759
rect 66103 67713 66181 67759
rect 66227 67713 66305 67759
rect 66351 67713 66429 67759
rect 66475 67713 66553 67759
rect 66599 67713 66677 67759
rect 66723 67713 66801 67759
rect 66847 67713 66925 67759
rect 66971 67713 67049 67759
rect 67095 67713 67173 67759
rect 67219 67713 67297 67759
rect 67343 67713 67421 67759
rect 67467 67713 67545 67759
rect 67591 67713 67669 67759
rect 67715 67713 67793 67759
rect 67839 67713 67917 67759
rect 67963 67713 68041 67759
rect 68087 67713 68165 67759
rect 68211 67713 68289 67759
rect 68335 67713 68413 67759
rect 68459 67713 68537 67759
rect 68583 67713 68661 67759
rect 68707 67713 68785 67759
rect 68831 67713 68909 67759
rect 68955 67713 69033 67759
rect 69079 67713 69157 67759
rect 69203 67713 69281 67759
rect 69327 67713 69405 67759
rect 69451 67713 69529 67759
rect 69575 67713 69653 67759
rect 69699 67713 69777 67759
rect 69823 67713 69901 67759
rect 69947 67713 70025 67759
rect 70071 67713 70149 67759
rect 70195 67713 70273 67759
rect 70319 67713 70397 67759
rect 70443 67713 70521 67759
rect 70567 67713 70645 67759
rect 70691 67713 70769 67759
rect 70815 67713 70893 67759
rect 70939 67713 71017 67759
rect 71063 67713 71141 67759
rect 71187 67713 71265 67759
rect 71311 67713 71389 67759
rect 71435 67713 71513 67759
rect 71559 67713 71637 67759
rect 71683 67713 71761 67759
rect 71807 67713 71885 67759
rect 71931 67713 72009 67759
rect 72055 67713 72133 67759
rect 72179 67713 72257 67759
rect 72303 67713 72381 67759
rect 72427 67713 72505 67759
rect 72551 67713 72629 67759
rect 72675 67713 72753 67759
rect 72799 67713 72877 67759
rect 72923 67713 73001 67759
rect 73047 67713 73125 67759
rect 73171 67713 73249 67759
rect 73295 67713 73373 67759
rect 73419 67713 73497 67759
rect 73543 67713 73621 67759
rect 73667 67713 73745 67759
rect 73791 67713 73869 67759
rect 73915 67713 73993 67759
rect 74039 67713 74117 67759
rect 74163 67713 74241 67759
rect 74287 67713 74365 67759
rect 74411 67713 74489 67759
rect 74535 67713 74613 67759
rect 74659 67713 74737 67759
rect 74783 67713 74861 67759
rect 74907 67713 74985 67759
rect 75031 67713 75109 67759
rect 75155 67713 75233 67759
rect 75279 67713 75357 67759
rect 75403 67713 75481 67759
rect 75527 67713 75605 67759
rect 75651 67713 75729 67759
rect 75775 67713 75853 67759
rect 75899 67713 75977 67759
rect 76023 67713 76101 67759
rect 76147 67713 76225 67759
rect 76271 67713 76349 67759
rect 76395 67713 76473 67759
rect 76519 67713 76597 67759
rect 76643 67713 76721 67759
rect 76767 67713 76845 67759
rect 76891 67713 76969 67759
rect 77015 67713 77093 67759
rect 77139 67713 77217 67759
rect 77263 67713 77341 67759
rect 77387 67713 77465 67759
rect 77511 67713 77589 67759
rect 77635 67713 77713 67759
rect 77759 67713 77837 67759
rect 77883 67713 77961 67759
rect 78007 67713 78085 67759
rect 78131 67713 78209 67759
rect 78255 67713 78333 67759
rect 78379 67713 78457 67759
rect 78503 67713 78581 67759
rect 78627 67713 78705 67759
rect 78751 67713 78829 67759
rect 78875 67713 78953 67759
rect 78999 67713 79077 67759
rect 79123 67713 79201 67759
rect 79247 67713 79325 67759
rect 79371 67713 79449 67759
rect 79495 67713 79573 67759
rect 79619 67713 79697 67759
rect 79743 67713 79821 67759
rect 79867 67713 79945 67759
rect 79991 67713 80069 67759
rect 80115 67713 80193 67759
rect 80239 67713 80317 67759
rect 80363 67713 80441 67759
rect 80487 67713 80565 67759
rect 80611 67713 80689 67759
rect 80735 67713 80813 67759
rect 80859 67713 80937 67759
rect 80983 67713 81061 67759
rect 81107 67713 81185 67759
rect 81231 67713 81309 67759
rect 81355 67713 81433 67759
rect 81479 67713 81557 67759
rect 81603 67713 81681 67759
rect 81727 67713 81805 67759
rect 81851 67713 81929 67759
rect 81975 67713 82053 67759
rect 82099 67713 82177 67759
rect 82223 67713 82301 67759
rect 82347 67713 82425 67759
rect 82471 67713 82549 67759
rect 82595 67713 82673 67759
rect 82719 67713 82797 67759
rect 82843 67713 82921 67759
rect 82967 67713 83045 67759
rect 83091 67713 83169 67759
rect 83215 67713 83293 67759
rect 83339 67713 83417 67759
rect 83463 67713 83541 67759
rect 83587 67713 83665 67759
rect 83711 67713 83789 67759
rect 83835 67713 83913 67759
rect 83959 67713 84037 67759
rect 84083 67713 84161 67759
rect 84207 67713 84285 67759
rect 84331 67713 84409 67759
rect 84455 67713 84533 67759
rect 84579 67713 84657 67759
rect 84703 67713 84781 67759
rect 84827 67713 84905 67759
rect 84951 67713 85029 67759
rect 85075 67713 85153 67759
rect 85199 67713 85277 67759
rect 85323 67713 85401 67759
rect 85447 67713 85525 67759
rect 85571 67713 85649 67759
rect 85695 67713 85808 67759
rect 0 67635 85808 67713
rect 0 67589 89 67635
rect 135 67589 213 67635
rect 259 67589 337 67635
rect 383 67589 461 67635
rect 507 67589 585 67635
rect 631 67589 709 67635
rect 755 67589 833 67635
rect 879 67589 957 67635
rect 1003 67589 1081 67635
rect 1127 67589 1205 67635
rect 1251 67589 1329 67635
rect 1375 67589 1453 67635
rect 1499 67589 1577 67635
rect 1623 67589 1701 67635
rect 1747 67589 1825 67635
rect 1871 67589 1949 67635
rect 1995 67589 2073 67635
rect 2119 67589 2197 67635
rect 2243 67589 2321 67635
rect 2367 67589 2445 67635
rect 2491 67589 2569 67635
rect 2615 67589 2693 67635
rect 2739 67589 2817 67635
rect 2863 67589 2941 67635
rect 2987 67589 3065 67635
rect 3111 67589 3189 67635
rect 3235 67589 3313 67635
rect 3359 67589 3437 67635
rect 3483 67589 3561 67635
rect 3607 67589 3685 67635
rect 3731 67589 3809 67635
rect 3855 67589 3933 67635
rect 3979 67589 4057 67635
rect 4103 67589 4181 67635
rect 4227 67589 4305 67635
rect 4351 67589 4429 67635
rect 4475 67589 4553 67635
rect 4599 67589 4677 67635
rect 4723 67589 4801 67635
rect 4847 67589 4925 67635
rect 4971 67589 5049 67635
rect 5095 67589 5173 67635
rect 5219 67589 5297 67635
rect 5343 67589 5421 67635
rect 5467 67589 5545 67635
rect 5591 67589 5669 67635
rect 5715 67589 5793 67635
rect 5839 67589 5917 67635
rect 5963 67589 6041 67635
rect 6087 67589 6165 67635
rect 6211 67589 6289 67635
rect 6335 67589 6413 67635
rect 6459 67589 6537 67635
rect 6583 67589 6661 67635
rect 6707 67589 6785 67635
rect 6831 67589 6909 67635
rect 6955 67589 7033 67635
rect 7079 67589 7157 67635
rect 7203 67589 7281 67635
rect 7327 67589 7405 67635
rect 7451 67589 7529 67635
rect 7575 67589 7653 67635
rect 7699 67589 7777 67635
rect 7823 67589 7901 67635
rect 7947 67589 8025 67635
rect 8071 67589 8149 67635
rect 8195 67589 8273 67635
rect 8319 67589 8397 67635
rect 8443 67589 8521 67635
rect 8567 67589 8645 67635
rect 8691 67589 8769 67635
rect 8815 67589 8893 67635
rect 8939 67589 9017 67635
rect 9063 67589 9141 67635
rect 9187 67589 9265 67635
rect 9311 67589 9389 67635
rect 9435 67589 9513 67635
rect 9559 67589 9637 67635
rect 9683 67589 9761 67635
rect 9807 67589 9885 67635
rect 9931 67589 10009 67635
rect 10055 67589 10133 67635
rect 10179 67589 10257 67635
rect 10303 67589 10381 67635
rect 10427 67589 10505 67635
rect 10551 67589 10629 67635
rect 10675 67589 10753 67635
rect 10799 67589 10877 67635
rect 10923 67589 11001 67635
rect 11047 67589 11125 67635
rect 11171 67589 11249 67635
rect 11295 67589 11373 67635
rect 11419 67589 11497 67635
rect 11543 67589 11621 67635
rect 11667 67589 11745 67635
rect 11791 67589 11869 67635
rect 11915 67589 11993 67635
rect 12039 67589 12117 67635
rect 12163 67589 12241 67635
rect 12287 67589 12365 67635
rect 12411 67589 12489 67635
rect 12535 67589 12613 67635
rect 12659 67589 12737 67635
rect 12783 67589 12861 67635
rect 12907 67589 12985 67635
rect 13031 67589 13109 67635
rect 13155 67589 13233 67635
rect 13279 67589 13357 67635
rect 13403 67589 13481 67635
rect 13527 67589 13605 67635
rect 13651 67589 13729 67635
rect 13775 67589 13853 67635
rect 13899 67589 13977 67635
rect 14023 67589 14101 67635
rect 14147 67589 14225 67635
rect 14271 67589 14349 67635
rect 14395 67589 14473 67635
rect 14519 67589 14597 67635
rect 14643 67589 14721 67635
rect 14767 67589 14845 67635
rect 14891 67589 14969 67635
rect 15015 67589 15093 67635
rect 15139 67589 15217 67635
rect 15263 67589 15341 67635
rect 15387 67589 15465 67635
rect 15511 67589 15589 67635
rect 15635 67589 15713 67635
rect 15759 67589 15837 67635
rect 15883 67589 15961 67635
rect 16007 67589 16085 67635
rect 16131 67589 16209 67635
rect 16255 67589 16333 67635
rect 16379 67589 16457 67635
rect 16503 67589 16581 67635
rect 16627 67589 16705 67635
rect 16751 67589 16829 67635
rect 16875 67589 16953 67635
rect 16999 67589 17077 67635
rect 17123 67589 17201 67635
rect 17247 67589 17325 67635
rect 17371 67589 17449 67635
rect 17495 67589 17573 67635
rect 17619 67589 17697 67635
rect 17743 67589 17821 67635
rect 17867 67589 17945 67635
rect 17991 67589 18069 67635
rect 18115 67589 18193 67635
rect 18239 67589 18317 67635
rect 18363 67589 18441 67635
rect 18487 67589 18565 67635
rect 18611 67589 18689 67635
rect 18735 67589 18813 67635
rect 18859 67589 18937 67635
rect 18983 67589 19061 67635
rect 19107 67589 19185 67635
rect 19231 67589 19309 67635
rect 19355 67589 19433 67635
rect 19479 67589 19557 67635
rect 19603 67589 19681 67635
rect 19727 67589 19805 67635
rect 19851 67589 19929 67635
rect 19975 67589 20053 67635
rect 20099 67589 20177 67635
rect 20223 67589 20301 67635
rect 20347 67589 20425 67635
rect 20471 67589 20549 67635
rect 20595 67589 20673 67635
rect 20719 67589 20797 67635
rect 20843 67589 20921 67635
rect 20967 67589 21045 67635
rect 21091 67589 21169 67635
rect 21215 67589 21293 67635
rect 21339 67589 21417 67635
rect 21463 67589 21541 67635
rect 21587 67589 21665 67635
rect 21711 67589 21789 67635
rect 21835 67589 21913 67635
rect 21959 67589 22037 67635
rect 22083 67589 22161 67635
rect 22207 67589 22285 67635
rect 22331 67589 22409 67635
rect 22455 67589 22533 67635
rect 22579 67589 22657 67635
rect 22703 67589 22781 67635
rect 22827 67589 22905 67635
rect 22951 67589 23029 67635
rect 23075 67589 23153 67635
rect 23199 67589 23277 67635
rect 23323 67589 23401 67635
rect 23447 67589 23525 67635
rect 23571 67589 23649 67635
rect 23695 67589 23773 67635
rect 23819 67589 23897 67635
rect 23943 67589 24021 67635
rect 24067 67589 24145 67635
rect 24191 67589 24269 67635
rect 24315 67589 24393 67635
rect 24439 67589 24517 67635
rect 24563 67589 24641 67635
rect 24687 67589 24765 67635
rect 24811 67589 24889 67635
rect 24935 67589 25013 67635
rect 25059 67589 25137 67635
rect 25183 67589 25261 67635
rect 25307 67589 25385 67635
rect 25431 67589 25509 67635
rect 25555 67589 25633 67635
rect 25679 67589 25757 67635
rect 25803 67589 25881 67635
rect 25927 67589 26005 67635
rect 26051 67589 26129 67635
rect 26175 67589 26253 67635
rect 26299 67589 26377 67635
rect 26423 67589 26501 67635
rect 26547 67589 26625 67635
rect 26671 67589 26749 67635
rect 26795 67589 26873 67635
rect 26919 67589 26997 67635
rect 27043 67589 27121 67635
rect 27167 67589 27245 67635
rect 27291 67589 27369 67635
rect 27415 67589 27493 67635
rect 27539 67589 27617 67635
rect 27663 67589 27741 67635
rect 27787 67589 27865 67635
rect 27911 67589 27989 67635
rect 28035 67589 28113 67635
rect 28159 67589 28237 67635
rect 28283 67589 28361 67635
rect 28407 67589 28485 67635
rect 28531 67589 28609 67635
rect 28655 67589 28733 67635
rect 28779 67589 28857 67635
rect 28903 67589 28981 67635
rect 29027 67589 29105 67635
rect 29151 67589 29229 67635
rect 29275 67589 29353 67635
rect 29399 67589 29477 67635
rect 29523 67589 29601 67635
rect 29647 67589 29725 67635
rect 29771 67589 29849 67635
rect 29895 67589 29973 67635
rect 30019 67589 30097 67635
rect 30143 67589 30221 67635
rect 30267 67589 30345 67635
rect 30391 67589 30469 67635
rect 30515 67589 30593 67635
rect 30639 67589 30717 67635
rect 30763 67589 30841 67635
rect 30887 67589 30965 67635
rect 31011 67589 31089 67635
rect 31135 67589 31213 67635
rect 31259 67589 31337 67635
rect 31383 67589 31461 67635
rect 31507 67589 31585 67635
rect 31631 67589 31709 67635
rect 31755 67589 31833 67635
rect 31879 67589 31957 67635
rect 32003 67589 32081 67635
rect 32127 67589 32205 67635
rect 32251 67589 32329 67635
rect 32375 67589 32453 67635
rect 32499 67589 32577 67635
rect 32623 67589 32701 67635
rect 32747 67589 32825 67635
rect 32871 67589 32949 67635
rect 32995 67589 33073 67635
rect 33119 67589 33197 67635
rect 33243 67589 33321 67635
rect 33367 67589 33445 67635
rect 33491 67589 33569 67635
rect 33615 67589 33693 67635
rect 33739 67589 33817 67635
rect 33863 67589 33941 67635
rect 33987 67589 34065 67635
rect 34111 67589 34189 67635
rect 34235 67589 34313 67635
rect 34359 67589 34437 67635
rect 34483 67589 34561 67635
rect 34607 67589 34685 67635
rect 34731 67589 34809 67635
rect 34855 67589 34933 67635
rect 34979 67589 35057 67635
rect 35103 67589 35181 67635
rect 35227 67589 35305 67635
rect 35351 67589 35429 67635
rect 35475 67589 35553 67635
rect 35599 67589 35677 67635
rect 35723 67589 35801 67635
rect 35847 67589 35925 67635
rect 35971 67589 36049 67635
rect 36095 67589 36173 67635
rect 36219 67589 36297 67635
rect 36343 67589 36421 67635
rect 36467 67589 36545 67635
rect 36591 67589 36669 67635
rect 36715 67589 36793 67635
rect 36839 67589 36917 67635
rect 36963 67589 37041 67635
rect 37087 67589 37165 67635
rect 37211 67589 37289 67635
rect 37335 67589 37413 67635
rect 37459 67589 37537 67635
rect 37583 67589 37661 67635
rect 37707 67589 37785 67635
rect 37831 67589 37909 67635
rect 37955 67589 38033 67635
rect 38079 67589 38157 67635
rect 38203 67589 38281 67635
rect 38327 67589 38405 67635
rect 38451 67589 38529 67635
rect 38575 67589 38653 67635
rect 38699 67589 38777 67635
rect 38823 67589 38901 67635
rect 38947 67589 39025 67635
rect 39071 67589 39149 67635
rect 39195 67589 39273 67635
rect 39319 67589 39397 67635
rect 39443 67589 39521 67635
rect 39567 67589 39645 67635
rect 39691 67589 39769 67635
rect 39815 67589 39893 67635
rect 39939 67589 40017 67635
rect 40063 67589 40141 67635
rect 40187 67589 40265 67635
rect 40311 67589 40389 67635
rect 40435 67589 40513 67635
rect 40559 67589 40637 67635
rect 40683 67589 40761 67635
rect 40807 67589 40885 67635
rect 40931 67589 41009 67635
rect 41055 67589 41133 67635
rect 41179 67589 41257 67635
rect 41303 67589 41381 67635
rect 41427 67589 41505 67635
rect 41551 67589 41629 67635
rect 41675 67589 41753 67635
rect 41799 67589 41877 67635
rect 41923 67589 42001 67635
rect 42047 67589 42125 67635
rect 42171 67589 42249 67635
rect 42295 67589 42373 67635
rect 42419 67589 42497 67635
rect 42543 67589 42621 67635
rect 42667 67589 42745 67635
rect 42791 67589 42869 67635
rect 42915 67589 42993 67635
rect 43039 67589 43117 67635
rect 43163 67589 43241 67635
rect 43287 67589 43365 67635
rect 43411 67589 43489 67635
rect 43535 67589 43613 67635
rect 43659 67589 43737 67635
rect 43783 67589 43861 67635
rect 43907 67589 43985 67635
rect 44031 67589 44109 67635
rect 44155 67589 44233 67635
rect 44279 67589 44357 67635
rect 44403 67589 44481 67635
rect 44527 67589 44605 67635
rect 44651 67589 44729 67635
rect 44775 67589 44853 67635
rect 44899 67589 44977 67635
rect 45023 67589 45101 67635
rect 45147 67589 45225 67635
rect 45271 67589 45349 67635
rect 45395 67589 45473 67635
rect 45519 67589 45597 67635
rect 45643 67589 45721 67635
rect 45767 67589 45845 67635
rect 45891 67589 45969 67635
rect 46015 67589 46093 67635
rect 46139 67589 46217 67635
rect 46263 67589 46341 67635
rect 46387 67589 46465 67635
rect 46511 67589 46589 67635
rect 46635 67589 46713 67635
rect 46759 67589 46837 67635
rect 46883 67589 46961 67635
rect 47007 67589 47085 67635
rect 47131 67589 47209 67635
rect 47255 67589 47333 67635
rect 47379 67589 47457 67635
rect 47503 67589 47581 67635
rect 47627 67589 47705 67635
rect 47751 67589 47829 67635
rect 47875 67589 47953 67635
rect 47999 67589 48077 67635
rect 48123 67589 48201 67635
rect 48247 67589 48325 67635
rect 48371 67589 48449 67635
rect 48495 67589 48573 67635
rect 48619 67589 48697 67635
rect 48743 67589 48821 67635
rect 48867 67589 48945 67635
rect 48991 67589 49069 67635
rect 49115 67589 49193 67635
rect 49239 67589 49317 67635
rect 49363 67589 49441 67635
rect 49487 67589 49565 67635
rect 49611 67589 49689 67635
rect 49735 67589 49813 67635
rect 49859 67589 49937 67635
rect 49983 67589 50061 67635
rect 50107 67589 50185 67635
rect 50231 67589 50309 67635
rect 50355 67589 50433 67635
rect 50479 67589 50557 67635
rect 50603 67589 50681 67635
rect 50727 67589 50805 67635
rect 50851 67589 50929 67635
rect 50975 67589 51053 67635
rect 51099 67589 51177 67635
rect 51223 67589 51301 67635
rect 51347 67589 51425 67635
rect 51471 67589 51549 67635
rect 51595 67589 51673 67635
rect 51719 67589 51797 67635
rect 51843 67589 51921 67635
rect 51967 67589 52045 67635
rect 52091 67589 52169 67635
rect 52215 67589 52293 67635
rect 52339 67589 52417 67635
rect 52463 67589 52541 67635
rect 52587 67589 52665 67635
rect 52711 67589 52789 67635
rect 52835 67589 52913 67635
rect 52959 67589 53037 67635
rect 53083 67589 53161 67635
rect 53207 67589 53285 67635
rect 53331 67589 53409 67635
rect 53455 67589 53533 67635
rect 53579 67589 53657 67635
rect 53703 67589 53781 67635
rect 53827 67589 53905 67635
rect 53951 67589 54029 67635
rect 54075 67589 54153 67635
rect 54199 67589 54277 67635
rect 54323 67589 54401 67635
rect 54447 67589 54525 67635
rect 54571 67589 54649 67635
rect 54695 67589 54773 67635
rect 54819 67589 54897 67635
rect 54943 67589 55021 67635
rect 55067 67589 55145 67635
rect 55191 67589 55269 67635
rect 55315 67589 55393 67635
rect 55439 67589 55517 67635
rect 55563 67589 55641 67635
rect 55687 67589 55765 67635
rect 55811 67589 55889 67635
rect 55935 67589 56013 67635
rect 56059 67589 56137 67635
rect 56183 67589 56261 67635
rect 56307 67589 56385 67635
rect 56431 67589 56509 67635
rect 56555 67589 56633 67635
rect 56679 67589 56757 67635
rect 56803 67589 56881 67635
rect 56927 67589 57005 67635
rect 57051 67589 57129 67635
rect 57175 67589 57253 67635
rect 57299 67589 57377 67635
rect 57423 67589 57501 67635
rect 57547 67589 57625 67635
rect 57671 67589 57749 67635
rect 57795 67589 57873 67635
rect 57919 67589 57997 67635
rect 58043 67589 58121 67635
rect 58167 67589 58245 67635
rect 58291 67589 58369 67635
rect 58415 67589 58493 67635
rect 58539 67589 58617 67635
rect 58663 67589 58741 67635
rect 58787 67589 58865 67635
rect 58911 67589 58989 67635
rect 59035 67589 59113 67635
rect 59159 67589 59237 67635
rect 59283 67589 59361 67635
rect 59407 67589 59485 67635
rect 59531 67589 59609 67635
rect 59655 67589 59733 67635
rect 59779 67589 59857 67635
rect 59903 67589 59981 67635
rect 60027 67589 60105 67635
rect 60151 67589 60229 67635
rect 60275 67589 60353 67635
rect 60399 67589 60477 67635
rect 60523 67589 60601 67635
rect 60647 67589 60725 67635
rect 60771 67589 60849 67635
rect 60895 67589 60973 67635
rect 61019 67589 61097 67635
rect 61143 67589 61221 67635
rect 61267 67589 61345 67635
rect 61391 67589 61469 67635
rect 61515 67589 61593 67635
rect 61639 67589 61717 67635
rect 61763 67589 61841 67635
rect 61887 67589 61965 67635
rect 62011 67589 62089 67635
rect 62135 67589 62213 67635
rect 62259 67589 62337 67635
rect 62383 67589 62461 67635
rect 62507 67589 62585 67635
rect 62631 67589 62709 67635
rect 62755 67589 62833 67635
rect 62879 67589 62957 67635
rect 63003 67589 63081 67635
rect 63127 67589 63205 67635
rect 63251 67589 63329 67635
rect 63375 67589 63453 67635
rect 63499 67589 63577 67635
rect 63623 67589 63701 67635
rect 63747 67589 63825 67635
rect 63871 67589 63949 67635
rect 63995 67589 64073 67635
rect 64119 67589 64197 67635
rect 64243 67589 64321 67635
rect 64367 67589 64445 67635
rect 64491 67589 64569 67635
rect 64615 67589 64693 67635
rect 64739 67589 64817 67635
rect 64863 67589 64941 67635
rect 64987 67589 65065 67635
rect 65111 67589 65189 67635
rect 65235 67589 65313 67635
rect 65359 67589 65437 67635
rect 65483 67589 65561 67635
rect 65607 67589 65685 67635
rect 65731 67589 65809 67635
rect 65855 67589 65933 67635
rect 65979 67589 66057 67635
rect 66103 67589 66181 67635
rect 66227 67589 66305 67635
rect 66351 67589 66429 67635
rect 66475 67589 66553 67635
rect 66599 67589 66677 67635
rect 66723 67589 66801 67635
rect 66847 67589 66925 67635
rect 66971 67589 67049 67635
rect 67095 67589 67173 67635
rect 67219 67589 67297 67635
rect 67343 67589 67421 67635
rect 67467 67589 67545 67635
rect 67591 67589 67669 67635
rect 67715 67589 67793 67635
rect 67839 67589 67917 67635
rect 67963 67589 68041 67635
rect 68087 67589 68165 67635
rect 68211 67589 68289 67635
rect 68335 67589 68413 67635
rect 68459 67589 68537 67635
rect 68583 67589 68661 67635
rect 68707 67589 68785 67635
rect 68831 67589 68909 67635
rect 68955 67589 69033 67635
rect 69079 67589 69157 67635
rect 69203 67589 69281 67635
rect 69327 67589 69405 67635
rect 69451 67589 69529 67635
rect 69575 67589 69653 67635
rect 69699 67589 69777 67635
rect 69823 67589 69901 67635
rect 69947 67589 70025 67635
rect 70071 67589 70149 67635
rect 70195 67589 70273 67635
rect 70319 67589 70397 67635
rect 70443 67589 70521 67635
rect 70567 67589 70645 67635
rect 70691 67589 70769 67635
rect 70815 67589 70893 67635
rect 70939 67589 71017 67635
rect 71063 67589 71141 67635
rect 71187 67589 71265 67635
rect 71311 67589 71389 67635
rect 71435 67589 71513 67635
rect 71559 67589 71637 67635
rect 71683 67589 71761 67635
rect 71807 67589 71885 67635
rect 71931 67589 72009 67635
rect 72055 67589 72133 67635
rect 72179 67589 72257 67635
rect 72303 67589 72381 67635
rect 72427 67589 72505 67635
rect 72551 67589 72629 67635
rect 72675 67589 72753 67635
rect 72799 67589 72877 67635
rect 72923 67589 73001 67635
rect 73047 67589 73125 67635
rect 73171 67589 73249 67635
rect 73295 67589 73373 67635
rect 73419 67589 73497 67635
rect 73543 67589 73621 67635
rect 73667 67589 73745 67635
rect 73791 67589 73869 67635
rect 73915 67589 73993 67635
rect 74039 67589 74117 67635
rect 74163 67589 74241 67635
rect 74287 67589 74365 67635
rect 74411 67589 74489 67635
rect 74535 67589 74613 67635
rect 74659 67589 74737 67635
rect 74783 67589 74861 67635
rect 74907 67589 74985 67635
rect 75031 67589 75109 67635
rect 75155 67589 75233 67635
rect 75279 67589 75357 67635
rect 75403 67589 75481 67635
rect 75527 67589 75605 67635
rect 75651 67589 75729 67635
rect 75775 67589 75853 67635
rect 75899 67589 75977 67635
rect 76023 67589 76101 67635
rect 76147 67589 76225 67635
rect 76271 67589 76349 67635
rect 76395 67589 76473 67635
rect 76519 67589 76597 67635
rect 76643 67589 76721 67635
rect 76767 67589 76845 67635
rect 76891 67589 76969 67635
rect 77015 67589 77093 67635
rect 77139 67589 77217 67635
rect 77263 67589 77341 67635
rect 77387 67589 77465 67635
rect 77511 67589 77589 67635
rect 77635 67589 77713 67635
rect 77759 67589 77837 67635
rect 77883 67589 77961 67635
rect 78007 67589 78085 67635
rect 78131 67589 78209 67635
rect 78255 67589 78333 67635
rect 78379 67589 78457 67635
rect 78503 67589 78581 67635
rect 78627 67589 78705 67635
rect 78751 67589 78829 67635
rect 78875 67589 78953 67635
rect 78999 67589 79077 67635
rect 79123 67589 79201 67635
rect 79247 67589 79325 67635
rect 79371 67589 79449 67635
rect 79495 67589 79573 67635
rect 79619 67589 79697 67635
rect 79743 67589 79821 67635
rect 79867 67589 79945 67635
rect 79991 67589 80069 67635
rect 80115 67589 80193 67635
rect 80239 67589 80317 67635
rect 80363 67589 80441 67635
rect 80487 67589 80565 67635
rect 80611 67589 80689 67635
rect 80735 67589 80813 67635
rect 80859 67589 80937 67635
rect 80983 67589 81061 67635
rect 81107 67589 81185 67635
rect 81231 67589 81309 67635
rect 81355 67589 81433 67635
rect 81479 67589 81557 67635
rect 81603 67589 81681 67635
rect 81727 67589 81805 67635
rect 81851 67589 81929 67635
rect 81975 67589 82053 67635
rect 82099 67589 82177 67635
rect 82223 67589 82301 67635
rect 82347 67589 82425 67635
rect 82471 67589 82549 67635
rect 82595 67589 82673 67635
rect 82719 67589 82797 67635
rect 82843 67589 82921 67635
rect 82967 67589 83045 67635
rect 83091 67589 83169 67635
rect 83215 67589 83293 67635
rect 83339 67589 83417 67635
rect 83463 67589 83541 67635
rect 83587 67589 83665 67635
rect 83711 67589 83789 67635
rect 83835 67589 83913 67635
rect 83959 67589 84037 67635
rect 84083 67589 84161 67635
rect 84207 67589 84285 67635
rect 84331 67589 84409 67635
rect 84455 67589 84533 67635
rect 84579 67589 84657 67635
rect 84703 67589 84781 67635
rect 84827 67589 84905 67635
rect 84951 67589 85029 67635
rect 85075 67589 85153 67635
rect 85199 67589 85277 67635
rect 85323 67589 85401 67635
rect 85447 67589 85525 67635
rect 85571 67589 85649 67635
rect 85695 67589 85808 67635
rect 0 67511 85808 67589
rect 0 67465 89 67511
rect 135 67465 213 67511
rect 259 67465 337 67511
rect 383 67465 461 67511
rect 507 67465 585 67511
rect 631 67465 709 67511
rect 755 67465 833 67511
rect 879 67465 957 67511
rect 1003 67465 1081 67511
rect 1127 67465 1205 67511
rect 1251 67465 1329 67511
rect 1375 67465 1453 67511
rect 1499 67465 1577 67511
rect 1623 67465 1701 67511
rect 1747 67465 1825 67511
rect 1871 67465 1949 67511
rect 1995 67465 2073 67511
rect 2119 67465 2197 67511
rect 2243 67465 2321 67511
rect 2367 67465 2445 67511
rect 2491 67465 2569 67511
rect 2615 67465 2693 67511
rect 2739 67465 2817 67511
rect 2863 67465 2941 67511
rect 2987 67465 3065 67511
rect 3111 67465 3189 67511
rect 3235 67465 3313 67511
rect 3359 67465 3437 67511
rect 3483 67465 3561 67511
rect 3607 67465 3685 67511
rect 3731 67465 3809 67511
rect 3855 67465 3933 67511
rect 3979 67465 4057 67511
rect 4103 67465 4181 67511
rect 4227 67465 4305 67511
rect 4351 67465 4429 67511
rect 4475 67465 4553 67511
rect 4599 67465 4677 67511
rect 4723 67465 4801 67511
rect 4847 67465 4925 67511
rect 4971 67465 5049 67511
rect 5095 67465 5173 67511
rect 5219 67465 5297 67511
rect 5343 67465 5421 67511
rect 5467 67465 5545 67511
rect 5591 67465 5669 67511
rect 5715 67465 5793 67511
rect 5839 67465 5917 67511
rect 5963 67465 6041 67511
rect 6087 67465 6165 67511
rect 6211 67465 6289 67511
rect 6335 67465 6413 67511
rect 6459 67465 6537 67511
rect 6583 67465 6661 67511
rect 6707 67465 6785 67511
rect 6831 67465 6909 67511
rect 6955 67465 7033 67511
rect 7079 67465 7157 67511
rect 7203 67465 7281 67511
rect 7327 67465 7405 67511
rect 7451 67465 7529 67511
rect 7575 67465 7653 67511
rect 7699 67465 7777 67511
rect 7823 67465 7901 67511
rect 7947 67465 8025 67511
rect 8071 67465 8149 67511
rect 8195 67465 8273 67511
rect 8319 67465 8397 67511
rect 8443 67465 8521 67511
rect 8567 67465 8645 67511
rect 8691 67465 8769 67511
rect 8815 67465 8893 67511
rect 8939 67465 9017 67511
rect 9063 67465 9141 67511
rect 9187 67465 9265 67511
rect 9311 67465 9389 67511
rect 9435 67465 9513 67511
rect 9559 67465 9637 67511
rect 9683 67465 9761 67511
rect 9807 67465 9885 67511
rect 9931 67465 10009 67511
rect 10055 67465 10133 67511
rect 10179 67465 10257 67511
rect 10303 67465 10381 67511
rect 10427 67465 10505 67511
rect 10551 67465 10629 67511
rect 10675 67465 10753 67511
rect 10799 67465 10877 67511
rect 10923 67465 11001 67511
rect 11047 67465 11125 67511
rect 11171 67465 11249 67511
rect 11295 67465 11373 67511
rect 11419 67465 11497 67511
rect 11543 67465 11621 67511
rect 11667 67465 11745 67511
rect 11791 67465 11869 67511
rect 11915 67465 11993 67511
rect 12039 67465 12117 67511
rect 12163 67465 12241 67511
rect 12287 67465 12365 67511
rect 12411 67465 12489 67511
rect 12535 67465 12613 67511
rect 12659 67465 12737 67511
rect 12783 67465 12861 67511
rect 12907 67465 12985 67511
rect 13031 67465 13109 67511
rect 13155 67465 13233 67511
rect 13279 67465 13357 67511
rect 13403 67465 13481 67511
rect 13527 67465 13605 67511
rect 13651 67465 13729 67511
rect 13775 67465 13853 67511
rect 13899 67465 13977 67511
rect 14023 67465 14101 67511
rect 14147 67465 14225 67511
rect 14271 67465 14349 67511
rect 14395 67465 14473 67511
rect 14519 67465 14597 67511
rect 14643 67465 14721 67511
rect 14767 67465 14845 67511
rect 14891 67465 14969 67511
rect 15015 67465 15093 67511
rect 15139 67465 15217 67511
rect 15263 67465 15341 67511
rect 15387 67465 15465 67511
rect 15511 67465 15589 67511
rect 15635 67465 15713 67511
rect 15759 67465 15837 67511
rect 15883 67465 15961 67511
rect 16007 67465 16085 67511
rect 16131 67465 16209 67511
rect 16255 67465 16333 67511
rect 16379 67465 16457 67511
rect 16503 67465 16581 67511
rect 16627 67465 16705 67511
rect 16751 67465 16829 67511
rect 16875 67465 16953 67511
rect 16999 67465 17077 67511
rect 17123 67465 17201 67511
rect 17247 67465 17325 67511
rect 17371 67465 17449 67511
rect 17495 67465 17573 67511
rect 17619 67465 17697 67511
rect 17743 67465 17821 67511
rect 17867 67465 17945 67511
rect 17991 67465 18069 67511
rect 18115 67465 18193 67511
rect 18239 67465 18317 67511
rect 18363 67465 18441 67511
rect 18487 67465 18565 67511
rect 18611 67465 18689 67511
rect 18735 67465 18813 67511
rect 18859 67465 18937 67511
rect 18983 67465 19061 67511
rect 19107 67465 19185 67511
rect 19231 67465 19309 67511
rect 19355 67465 19433 67511
rect 19479 67465 19557 67511
rect 19603 67465 19681 67511
rect 19727 67465 19805 67511
rect 19851 67465 19929 67511
rect 19975 67465 20053 67511
rect 20099 67465 20177 67511
rect 20223 67465 20301 67511
rect 20347 67465 20425 67511
rect 20471 67465 20549 67511
rect 20595 67465 20673 67511
rect 20719 67465 20797 67511
rect 20843 67465 20921 67511
rect 20967 67465 21045 67511
rect 21091 67465 21169 67511
rect 21215 67465 21293 67511
rect 21339 67465 21417 67511
rect 21463 67465 21541 67511
rect 21587 67465 21665 67511
rect 21711 67465 21789 67511
rect 21835 67465 21913 67511
rect 21959 67465 22037 67511
rect 22083 67465 22161 67511
rect 22207 67465 22285 67511
rect 22331 67465 22409 67511
rect 22455 67465 22533 67511
rect 22579 67465 22657 67511
rect 22703 67465 22781 67511
rect 22827 67465 22905 67511
rect 22951 67465 23029 67511
rect 23075 67465 23153 67511
rect 23199 67465 23277 67511
rect 23323 67465 23401 67511
rect 23447 67465 23525 67511
rect 23571 67465 23649 67511
rect 23695 67465 23773 67511
rect 23819 67465 23897 67511
rect 23943 67465 24021 67511
rect 24067 67465 24145 67511
rect 24191 67465 24269 67511
rect 24315 67465 24393 67511
rect 24439 67465 24517 67511
rect 24563 67465 24641 67511
rect 24687 67465 24765 67511
rect 24811 67465 24889 67511
rect 24935 67465 25013 67511
rect 25059 67465 25137 67511
rect 25183 67465 25261 67511
rect 25307 67465 25385 67511
rect 25431 67465 25509 67511
rect 25555 67465 25633 67511
rect 25679 67465 25757 67511
rect 25803 67465 25881 67511
rect 25927 67465 26005 67511
rect 26051 67465 26129 67511
rect 26175 67465 26253 67511
rect 26299 67465 26377 67511
rect 26423 67465 26501 67511
rect 26547 67465 26625 67511
rect 26671 67465 26749 67511
rect 26795 67465 26873 67511
rect 26919 67465 26997 67511
rect 27043 67465 27121 67511
rect 27167 67465 27245 67511
rect 27291 67465 27369 67511
rect 27415 67465 27493 67511
rect 27539 67465 27617 67511
rect 27663 67465 27741 67511
rect 27787 67465 27865 67511
rect 27911 67465 27989 67511
rect 28035 67465 28113 67511
rect 28159 67465 28237 67511
rect 28283 67465 28361 67511
rect 28407 67465 28485 67511
rect 28531 67465 28609 67511
rect 28655 67465 28733 67511
rect 28779 67465 28857 67511
rect 28903 67465 28981 67511
rect 29027 67465 29105 67511
rect 29151 67465 29229 67511
rect 29275 67465 29353 67511
rect 29399 67465 29477 67511
rect 29523 67465 29601 67511
rect 29647 67465 29725 67511
rect 29771 67465 29849 67511
rect 29895 67465 29973 67511
rect 30019 67465 30097 67511
rect 30143 67465 30221 67511
rect 30267 67465 30345 67511
rect 30391 67465 30469 67511
rect 30515 67465 30593 67511
rect 30639 67465 30717 67511
rect 30763 67465 30841 67511
rect 30887 67465 30965 67511
rect 31011 67465 31089 67511
rect 31135 67465 31213 67511
rect 31259 67465 31337 67511
rect 31383 67465 31461 67511
rect 31507 67465 31585 67511
rect 31631 67465 31709 67511
rect 31755 67465 31833 67511
rect 31879 67465 31957 67511
rect 32003 67465 32081 67511
rect 32127 67465 32205 67511
rect 32251 67465 32329 67511
rect 32375 67465 32453 67511
rect 32499 67465 32577 67511
rect 32623 67465 32701 67511
rect 32747 67465 32825 67511
rect 32871 67465 32949 67511
rect 32995 67465 33073 67511
rect 33119 67465 33197 67511
rect 33243 67465 33321 67511
rect 33367 67465 33445 67511
rect 33491 67465 33569 67511
rect 33615 67465 33693 67511
rect 33739 67465 33817 67511
rect 33863 67465 33941 67511
rect 33987 67465 34065 67511
rect 34111 67465 34189 67511
rect 34235 67465 34313 67511
rect 34359 67465 34437 67511
rect 34483 67465 34561 67511
rect 34607 67465 34685 67511
rect 34731 67465 34809 67511
rect 34855 67465 34933 67511
rect 34979 67465 35057 67511
rect 35103 67465 35181 67511
rect 35227 67465 35305 67511
rect 35351 67465 35429 67511
rect 35475 67465 35553 67511
rect 35599 67465 35677 67511
rect 35723 67465 35801 67511
rect 35847 67465 35925 67511
rect 35971 67465 36049 67511
rect 36095 67465 36173 67511
rect 36219 67465 36297 67511
rect 36343 67465 36421 67511
rect 36467 67465 36545 67511
rect 36591 67465 36669 67511
rect 36715 67465 36793 67511
rect 36839 67465 36917 67511
rect 36963 67465 37041 67511
rect 37087 67465 37165 67511
rect 37211 67465 37289 67511
rect 37335 67465 37413 67511
rect 37459 67465 37537 67511
rect 37583 67465 37661 67511
rect 37707 67465 37785 67511
rect 37831 67465 37909 67511
rect 37955 67465 38033 67511
rect 38079 67465 38157 67511
rect 38203 67465 38281 67511
rect 38327 67465 38405 67511
rect 38451 67465 38529 67511
rect 38575 67465 38653 67511
rect 38699 67465 38777 67511
rect 38823 67465 38901 67511
rect 38947 67465 39025 67511
rect 39071 67465 39149 67511
rect 39195 67465 39273 67511
rect 39319 67465 39397 67511
rect 39443 67465 39521 67511
rect 39567 67465 39645 67511
rect 39691 67465 39769 67511
rect 39815 67465 39893 67511
rect 39939 67465 40017 67511
rect 40063 67465 40141 67511
rect 40187 67465 40265 67511
rect 40311 67465 40389 67511
rect 40435 67465 40513 67511
rect 40559 67465 40637 67511
rect 40683 67465 40761 67511
rect 40807 67465 40885 67511
rect 40931 67465 41009 67511
rect 41055 67465 41133 67511
rect 41179 67465 41257 67511
rect 41303 67465 41381 67511
rect 41427 67465 41505 67511
rect 41551 67465 41629 67511
rect 41675 67465 41753 67511
rect 41799 67465 41877 67511
rect 41923 67465 42001 67511
rect 42047 67465 42125 67511
rect 42171 67465 42249 67511
rect 42295 67465 42373 67511
rect 42419 67465 42497 67511
rect 42543 67465 42621 67511
rect 42667 67465 42745 67511
rect 42791 67465 42869 67511
rect 42915 67465 42993 67511
rect 43039 67465 43117 67511
rect 43163 67465 43241 67511
rect 43287 67465 43365 67511
rect 43411 67465 43489 67511
rect 43535 67465 43613 67511
rect 43659 67465 43737 67511
rect 43783 67465 43861 67511
rect 43907 67465 43985 67511
rect 44031 67465 44109 67511
rect 44155 67465 44233 67511
rect 44279 67465 44357 67511
rect 44403 67465 44481 67511
rect 44527 67465 44605 67511
rect 44651 67465 44729 67511
rect 44775 67465 44853 67511
rect 44899 67465 44977 67511
rect 45023 67465 45101 67511
rect 45147 67465 45225 67511
rect 45271 67465 45349 67511
rect 45395 67465 45473 67511
rect 45519 67465 45597 67511
rect 45643 67465 45721 67511
rect 45767 67465 45845 67511
rect 45891 67465 45969 67511
rect 46015 67465 46093 67511
rect 46139 67465 46217 67511
rect 46263 67465 46341 67511
rect 46387 67465 46465 67511
rect 46511 67465 46589 67511
rect 46635 67465 46713 67511
rect 46759 67465 46837 67511
rect 46883 67465 46961 67511
rect 47007 67465 47085 67511
rect 47131 67465 47209 67511
rect 47255 67465 47333 67511
rect 47379 67465 47457 67511
rect 47503 67465 47581 67511
rect 47627 67465 47705 67511
rect 47751 67465 47829 67511
rect 47875 67465 47953 67511
rect 47999 67465 48077 67511
rect 48123 67465 48201 67511
rect 48247 67465 48325 67511
rect 48371 67465 48449 67511
rect 48495 67465 48573 67511
rect 48619 67465 48697 67511
rect 48743 67465 48821 67511
rect 48867 67465 48945 67511
rect 48991 67465 49069 67511
rect 49115 67465 49193 67511
rect 49239 67465 49317 67511
rect 49363 67465 49441 67511
rect 49487 67465 49565 67511
rect 49611 67465 49689 67511
rect 49735 67465 49813 67511
rect 49859 67465 49937 67511
rect 49983 67465 50061 67511
rect 50107 67465 50185 67511
rect 50231 67465 50309 67511
rect 50355 67465 50433 67511
rect 50479 67465 50557 67511
rect 50603 67465 50681 67511
rect 50727 67465 50805 67511
rect 50851 67465 50929 67511
rect 50975 67465 51053 67511
rect 51099 67465 51177 67511
rect 51223 67465 51301 67511
rect 51347 67465 51425 67511
rect 51471 67465 51549 67511
rect 51595 67465 51673 67511
rect 51719 67465 51797 67511
rect 51843 67465 51921 67511
rect 51967 67465 52045 67511
rect 52091 67465 52169 67511
rect 52215 67465 52293 67511
rect 52339 67465 52417 67511
rect 52463 67465 52541 67511
rect 52587 67465 52665 67511
rect 52711 67465 52789 67511
rect 52835 67465 52913 67511
rect 52959 67465 53037 67511
rect 53083 67465 53161 67511
rect 53207 67465 53285 67511
rect 53331 67465 53409 67511
rect 53455 67465 53533 67511
rect 53579 67465 53657 67511
rect 53703 67465 53781 67511
rect 53827 67465 53905 67511
rect 53951 67465 54029 67511
rect 54075 67465 54153 67511
rect 54199 67465 54277 67511
rect 54323 67465 54401 67511
rect 54447 67465 54525 67511
rect 54571 67465 54649 67511
rect 54695 67465 54773 67511
rect 54819 67465 54897 67511
rect 54943 67465 55021 67511
rect 55067 67465 55145 67511
rect 55191 67465 55269 67511
rect 55315 67465 55393 67511
rect 55439 67465 55517 67511
rect 55563 67465 55641 67511
rect 55687 67465 55765 67511
rect 55811 67465 55889 67511
rect 55935 67465 56013 67511
rect 56059 67465 56137 67511
rect 56183 67465 56261 67511
rect 56307 67465 56385 67511
rect 56431 67465 56509 67511
rect 56555 67465 56633 67511
rect 56679 67465 56757 67511
rect 56803 67465 56881 67511
rect 56927 67465 57005 67511
rect 57051 67465 57129 67511
rect 57175 67465 57253 67511
rect 57299 67465 57377 67511
rect 57423 67465 57501 67511
rect 57547 67465 57625 67511
rect 57671 67465 57749 67511
rect 57795 67465 57873 67511
rect 57919 67465 57997 67511
rect 58043 67465 58121 67511
rect 58167 67465 58245 67511
rect 58291 67465 58369 67511
rect 58415 67465 58493 67511
rect 58539 67465 58617 67511
rect 58663 67465 58741 67511
rect 58787 67465 58865 67511
rect 58911 67465 58989 67511
rect 59035 67465 59113 67511
rect 59159 67465 59237 67511
rect 59283 67465 59361 67511
rect 59407 67465 59485 67511
rect 59531 67465 59609 67511
rect 59655 67465 59733 67511
rect 59779 67465 59857 67511
rect 59903 67465 59981 67511
rect 60027 67465 60105 67511
rect 60151 67465 60229 67511
rect 60275 67465 60353 67511
rect 60399 67465 60477 67511
rect 60523 67465 60601 67511
rect 60647 67465 60725 67511
rect 60771 67465 60849 67511
rect 60895 67465 60973 67511
rect 61019 67465 61097 67511
rect 61143 67465 61221 67511
rect 61267 67465 61345 67511
rect 61391 67465 61469 67511
rect 61515 67465 61593 67511
rect 61639 67465 61717 67511
rect 61763 67465 61841 67511
rect 61887 67465 61965 67511
rect 62011 67465 62089 67511
rect 62135 67465 62213 67511
rect 62259 67465 62337 67511
rect 62383 67465 62461 67511
rect 62507 67465 62585 67511
rect 62631 67465 62709 67511
rect 62755 67465 62833 67511
rect 62879 67465 62957 67511
rect 63003 67465 63081 67511
rect 63127 67465 63205 67511
rect 63251 67465 63329 67511
rect 63375 67465 63453 67511
rect 63499 67465 63577 67511
rect 63623 67465 63701 67511
rect 63747 67465 63825 67511
rect 63871 67465 63949 67511
rect 63995 67465 64073 67511
rect 64119 67465 64197 67511
rect 64243 67465 64321 67511
rect 64367 67465 64445 67511
rect 64491 67465 64569 67511
rect 64615 67465 64693 67511
rect 64739 67465 64817 67511
rect 64863 67465 64941 67511
rect 64987 67465 65065 67511
rect 65111 67465 65189 67511
rect 65235 67465 65313 67511
rect 65359 67465 65437 67511
rect 65483 67465 65561 67511
rect 65607 67465 65685 67511
rect 65731 67465 65809 67511
rect 65855 67465 65933 67511
rect 65979 67465 66057 67511
rect 66103 67465 66181 67511
rect 66227 67465 66305 67511
rect 66351 67465 66429 67511
rect 66475 67465 66553 67511
rect 66599 67465 66677 67511
rect 66723 67465 66801 67511
rect 66847 67465 66925 67511
rect 66971 67465 67049 67511
rect 67095 67465 67173 67511
rect 67219 67465 67297 67511
rect 67343 67465 67421 67511
rect 67467 67465 67545 67511
rect 67591 67465 67669 67511
rect 67715 67465 67793 67511
rect 67839 67465 67917 67511
rect 67963 67465 68041 67511
rect 68087 67465 68165 67511
rect 68211 67465 68289 67511
rect 68335 67465 68413 67511
rect 68459 67465 68537 67511
rect 68583 67465 68661 67511
rect 68707 67465 68785 67511
rect 68831 67465 68909 67511
rect 68955 67465 69033 67511
rect 69079 67465 69157 67511
rect 69203 67465 69281 67511
rect 69327 67465 69405 67511
rect 69451 67465 69529 67511
rect 69575 67465 69653 67511
rect 69699 67465 69777 67511
rect 69823 67465 69901 67511
rect 69947 67465 70025 67511
rect 70071 67465 70149 67511
rect 70195 67465 70273 67511
rect 70319 67465 70397 67511
rect 70443 67465 70521 67511
rect 70567 67465 70645 67511
rect 70691 67465 70769 67511
rect 70815 67465 70893 67511
rect 70939 67465 71017 67511
rect 71063 67465 71141 67511
rect 71187 67465 71265 67511
rect 71311 67465 71389 67511
rect 71435 67465 71513 67511
rect 71559 67465 71637 67511
rect 71683 67465 71761 67511
rect 71807 67465 71885 67511
rect 71931 67465 72009 67511
rect 72055 67465 72133 67511
rect 72179 67465 72257 67511
rect 72303 67465 72381 67511
rect 72427 67465 72505 67511
rect 72551 67465 72629 67511
rect 72675 67465 72753 67511
rect 72799 67465 72877 67511
rect 72923 67465 73001 67511
rect 73047 67465 73125 67511
rect 73171 67465 73249 67511
rect 73295 67465 73373 67511
rect 73419 67465 73497 67511
rect 73543 67465 73621 67511
rect 73667 67465 73745 67511
rect 73791 67465 73869 67511
rect 73915 67465 73993 67511
rect 74039 67465 74117 67511
rect 74163 67465 74241 67511
rect 74287 67465 74365 67511
rect 74411 67465 74489 67511
rect 74535 67465 74613 67511
rect 74659 67465 74737 67511
rect 74783 67465 74861 67511
rect 74907 67465 74985 67511
rect 75031 67465 75109 67511
rect 75155 67465 75233 67511
rect 75279 67465 75357 67511
rect 75403 67465 75481 67511
rect 75527 67465 75605 67511
rect 75651 67465 75729 67511
rect 75775 67465 75853 67511
rect 75899 67465 75977 67511
rect 76023 67465 76101 67511
rect 76147 67465 76225 67511
rect 76271 67465 76349 67511
rect 76395 67465 76473 67511
rect 76519 67465 76597 67511
rect 76643 67465 76721 67511
rect 76767 67465 76845 67511
rect 76891 67465 76969 67511
rect 77015 67465 77093 67511
rect 77139 67465 77217 67511
rect 77263 67465 77341 67511
rect 77387 67465 77465 67511
rect 77511 67465 77589 67511
rect 77635 67465 77713 67511
rect 77759 67465 77837 67511
rect 77883 67465 77961 67511
rect 78007 67465 78085 67511
rect 78131 67465 78209 67511
rect 78255 67465 78333 67511
rect 78379 67465 78457 67511
rect 78503 67465 78581 67511
rect 78627 67465 78705 67511
rect 78751 67465 78829 67511
rect 78875 67465 78953 67511
rect 78999 67465 79077 67511
rect 79123 67465 79201 67511
rect 79247 67465 79325 67511
rect 79371 67465 79449 67511
rect 79495 67465 79573 67511
rect 79619 67465 79697 67511
rect 79743 67465 79821 67511
rect 79867 67465 79945 67511
rect 79991 67465 80069 67511
rect 80115 67465 80193 67511
rect 80239 67465 80317 67511
rect 80363 67465 80441 67511
rect 80487 67465 80565 67511
rect 80611 67465 80689 67511
rect 80735 67465 80813 67511
rect 80859 67465 80937 67511
rect 80983 67465 81061 67511
rect 81107 67465 81185 67511
rect 81231 67465 81309 67511
rect 81355 67465 81433 67511
rect 81479 67465 81557 67511
rect 81603 67465 81681 67511
rect 81727 67465 81805 67511
rect 81851 67465 81929 67511
rect 81975 67465 82053 67511
rect 82099 67465 82177 67511
rect 82223 67465 82301 67511
rect 82347 67465 82425 67511
rect 82471 67465 82549 67511
rect 82595 67465 82673 67511
rect 82719 67465 82797 67511
rect 82843 67465 82921 67511
rect 82967 67465 83045 67511
rect 83091 67465 83169 67511
rect 83215 67465 83293 67511
rect 83339 67465 83417 67511
rect 83463 67465 83541 67511
rect 83587 67465 83665 67511
rect 83711 67465 83789 67511
rect 83835 67465 83913 67511
rect 83959 67465 84037 67511
rect 84083 67465 84161 67511
rect 84207 67465 84285 67511
rect 84331 67465 84409 67511
rect 84455 67465 84533 67511
rect 84579 67465 84657 67511
rect 84703 67465 84781 67511
rect 84827 67465 84905 67511
rect 84951 67465 85029 67511
rect 85075 67465 85153 67511
rect 85199 67465 85277 67511
rect 85323 67465 85401 67511
rect 85447 67465 85525 67511
rect 85571 67465 85649 67511
rect 85695 67465 85808 67511
rect 0 67454 85808 67465
rect 0 67363 1000 67454
rect 0 1117 89 67363
rect 435 1117 1000 67363
rect 0 1026 1000 1117
rect 27105 67363 27473 67374
rect 27105 1117 27116 67363
rect 27462 1117 27473 67363
rect 57013 67363 57381 67374
rect 27553 67342 28421 67353
rect 27553 35996 27564 67342
rect 28410 35996 28421 67342
rect 27553 35985 28421 35996
rect 56099 67342 56967 67353
rect 56099 35996 56110 67342
rect 56956 35996 56967 67342
rect 56099 35985 56967 35996
rect 27553 34588 56921 34599
rect 27553 34242 27564 34588
rect 56910 34242 56921 34588
rect 27553 34231 56921 34242
rect 27105 1106 27473 1117
rect 57013 1117 57024 67363
rect 57370 1117 57381 67363
rect 57013 1106 57381 1117
rect 84808 67363 85808 67454
rect 84808 1117 85451 67363
rect 85797 1117 85808 67363
rect 84808 1026 85808 1117
rect 0 1015 85808 1026
rect 0 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85808 1015
rect 0 891 85808 969
rect 0 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85808 891
rect 0 767 85808 845
rect 0 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85808 767
rect 0 643 85808 721
rect 0 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85808 643
rect 0 586 85808 597
rect 0 403 1000 586
rect 84808 403 85808 586
<< metal2 >>
rect 424 403 1424 67376
rect 84384 403 85384 67376
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_0
timestamp 1755724134
transform 1 0 85474 0 1 1140
box 0 0 1 1
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_1
timestamp 1755724134
transform 1 0 27139 0 1 1140
box 0 0 1 1
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_2
timestamp 1755724134
transform 1 0 57047 0 1 1140
box 0 0 1 1
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_3
timestamp 1755724134
transform 1 0 112 0 1 1140
box 0 0 1 1
use M1_PSUB43105908781106_256x8m81  M1_PSUB43105908781106_256x8m81_0
timestamp 1755724134
transform 1 0 27587 0 1 34265
box 0 0 1 1
use M1_PSUB43105908781107_256x8m81  M1_PSUB43105908781107_256x8m81_0
timestamp 1755724134
transform 1 0 56133 0 1 36019
box 0 0 1 1
use M1_PSUB43105908781107_256x8m81  M1_PSUB43105908781107_256x8m81_1
timestamp 1755724134
transform 1 0 27587 0 1 36019
box 0 0 1 1
use M1_PSUB43105908781108_256x8m81  M1_PSUB43105908781108_256x8m81_0
timestamp 1755724134
transform 1 0 112 0 1 67488
box 0 0 1 1
use M1_PSUB43105908781108_256x8m81  M1_PSUB43105908781108_256x8m81_1
timestamp 1755724134
transform 1 0 112 0 1 620
box 0 0 1 1
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 448 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2141372
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2140118
string path 4.620 11.160 4.620 0.000 
<< end >>
