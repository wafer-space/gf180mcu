magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nbase >>
rect -1180 -1180 1180 1180
<< pdiff >>
rect -1000 973 1000 1000
rect -1000 -973 -973 973
rect 973 -973 1000 973
rect -1000 -1000 1000 -973
<< pdiffc >>
rect -973 -973 973 973
<< psubdiff >>
rect -1296 1277 1296 1296
rect -1296 1245 -1151 1277
rect -1296 -1245 -1277 1245
rect -1231 1231 -1151 1245
rect 1151 1245 1296 1277
rect 1151 1231 1231 1245
rect -1231 1212 1231 1231
rect -1231 -1212 -1212 1212
rect 1212 -1212 1231 1212
rect -1231 -1231 1231 -1212
rect -1231 -1245 -1151 -1231
rect -1296 -1277 -1151 -1245
rect 1151 -1245 1231 -1231
rect 1277 -1245 1296 1245
rect 1151 -1277 1296 -1245
rect -1296 -1296 1296 -1277
<< nsubdiff >>
rect -1148 1129 1148 1148
rect -1148 1104 -963 1129
rect -1148 -1104 -1129 1104
rect -1083 1083 -963 1104
rect 963 1104 1148 1129
rect 963 1083 1083 1104
rect -1083 1064 1083 1083
rect -1083 -1064 -1064 1064
rect 1064 -1064 1083 1064
rect -1083 -1083 1083 -1064
rect -1083 -1104 -963 -1083
rect -1148 -1129 -963 -1104
rect 963 -1104 1083 -1083
rect 1129 -1104 1148 1104
rect 963 -1129 1148 -1104
rect -1148 -1148 1148 -1129
<< psubdiffcont >>
rect -1277 -1245 -1231 1245
rect -1151 1231 1151 1277
rect -1151 -1277 1151 -1231
rect 1231 -1245 1277 1245
<< nsubdiffcont >>
rect -1129 -1104 -1083 1104
rect -963 1083 963 1129
rect -963 -1129 963 -1083
rect 1083 -1104 1129 1104
<< metal1 >>
rect -1296 1277 1296 1296
rect -1296 1245 -1151 1277
rect -1296 -1245 -1277 1245
rect -1231 1231 -1151 1245
rect 1151 1245 1296 1277
rect 1151 1231 1231 1245
rect -1231 1212 1231 1231
rect -1231 -1212 -1212 1212
rect -1148 1129 1148 1148
rect -1148 1104 -963 1129
rect -1148 -1104 -1129 1104
rect -1083 1083 -963 1104
rect 963 1104 1148 1129
rect 963 1083 1083 1104
rect -1083 1064 1083 1083
rect -1083 -1064 -1064 1064
rect -1000 973 1000 1000
rect -1000 -973 -973 973
rect 973 -973 1000 973
rect -1000 -1000 1000 -973
rect 1064 -1064 1083 1064
rect -1083 -1083 1083 -1064
rect -1083 -1104 -963 -1083
rect -1148 -1129 -963 -1104
rect 963 -1104 1083 -1083
rect 1129 -1104 1148 1104
rect 963 -1129 1148 -1104
rect -1148 -1148 1148 -1129
rect 1212 -1212 1231 1212
rect -1231 -1231 1231 -1212
rect -1231 -1245 -1151 -1231
rect -1296 -1277 -1151 -1245
rect 1151 -1245 1231 -1231
rect 1277 -1245 1296 1245
rect 1151 -1277 1296 -1245
rect -1296 -1296 1296 -1277
<< labels >>
flabel pdiffc 0 2 0 2 0 FreeSans 400 0 0 0 E
flabel nsubdiffcont 5 1113 5 1113 0 FreeSans 400 0 0 0 B
flabel nsubdiffcont 1106 2 1106 2 0 FreeSans 400 0 0 0 B
flabel nsubdiffcont -15 -1109 -15 -1109 0 FreeSans 400 0 0 0 B
flabel nsubdiffcont -1101 -2 -1101 -2 0 FreeSans 400 0 0 0 B
flabel psubdiffcont -5 1260 -5 1260 0 FreeSans 400 0 0 0 C
flabel psubdiffcont 1258 2 1258 2 0 FreeSans 400 0 0 0 C
flabel psubdiffcont 0 -1260 0 -1260 0 FreeSans 400 0 0 0 C
flabel psubdiffcont -1263 7 -1263 7 0 FreeSans 400 0 0 0 C
<< properties >>
string GDS_END 40322
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/pnp_10p00x10p00.gds
string GDS_START 112
string gencell pnp_10p00x10p00
string library gf180mcu
string parameter m=1
<< end >>
