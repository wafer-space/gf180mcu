magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
<< nwell >>
rect -86 355 3894 870
rect -86 352 952 355
rect 1550 352 3894 355
<< pwell >>
rect 952 352 1550 355
rect -86 -86 3894 352
<< mvnmos >>
rect 124 137 244 216
rect 348 137 468 216
rect 572 137 692 216
rect 799 137 919 216
rect 1059 156 1179 235
rect 1315 156 1435 235
rect 1815 91 1935 170
rect 2039 91 2159 170
rect 2407 91 2527 217
rect 2591 91 2711 217
rect 2815 91 2935 217
rect 3039 91 3159 217
rect 3263 91 3383 217
rect 3487 91 3607 217
<< mvpmos >>
rect 144 475 244 660
rect 348 475 448 660
rect 588 507 688 660
rect 887 507 987 660
rect 1127 475 1227 628
rect 1335 475 1435 628
rect 1809 475 1909 659
rect 2014 475 2114 659
rect 2407 472 2507 716
rect 2611 472 2711 716
rect 2815 472 2915 716
rect 3019 472 3119 716
rect 3223 472 3323 716
rect 3427 472 3527 716
<< mvndiff >>
rect 979 216 1059 235
rect 36 199 124 216
rect 36 153 49 199
rect 95 153 124 199
rect 36 137 124 153
rect 244 199 348 216
rect 244 153 273 199
rect 319 153 348 199
rect 244 137 348 153
rect 468 199 572 216
rect 468 153 497 199
rect 543 153 572 199
rect 468 137 572 153
rect 692 199 799 216
rect 692 153 721 199
rect 767 153 799 199
rect 692 137 799 153
rect 919 156 1059 216
rect 1179 215 1315 235
rect 1179 169 1224 215
rect 1270 169 1315 215
rect 1179 156 1315 169
rect 1435 215 1523 235
rect 1435 169 1464 215
rect 1510 169 1523 215
rect 1435 156 1523 169
rect 919 137 999 156
rect 1727 152 1815 170
rect 1727 106 1740 152
rect 1786 106 1815 152
rect 1727 91 1815 106
rect 1935 152 2039 170
rect 1935 106 1964 152
rect 2010 106 2039 152
rect 1935 91 2039 106
rect 2159 152 2247 170
rect 2159 106 2188 152
rect 2234 106 2247 152
rect 2159 91 2247 106
rect 2319 152 2407 217
rect 2319 106 2332 152
rect 2378 106 2407 152
rect 2319 91 2407 106
rect 2527 91 2591 217
rect 2711 150 2815 217
rect 2711 104 2740 150
rect 2786 104 2815 150
rect 2711 91 2815 104
rect 2935 198 3039 217
rect 2935 152 2964 198
rect 3010 152 3039 198
rect 2935 91 3039 152
rect 3159 150 3263 217
rect 3159 104 3188 150
rect 3234 104 3263 150
rect 3159 91 3263 104
rect 3383 198 3487 217
rect 3383 152 3412 198
rect 3458 152 3487 198
rect 3383 91 3487 152
rect 3607 150 3695 217
rect 3607 104 3636 150
rect 3682 104 3695 150
rect 3607 91 3695 104
<< mvpdiff >>
rect 56 647 144 660
rect 56 507 69 647
rect 115 507 144 647
rect 56 475 144 507
rect 244 475 348 660
rect 448 507 588 660
rect 688 614 887 660
rect 688 568 762 614
rect 808 568 887 614
rect 688 507 887 568
rect 987 628 1067 660
rect 2314 703 2407 716
rect 987 507 1127 628
rect 448 475 528 507
rect 1047 475 1127 507
rect 1227 578 1335 628
rect 1227 532 1256 578
rect 1302 532 1335 578
rect 1227 475 1335 532
rect 1435 544 1523 628
rect 1435 498 1464 544
rect 1510 498 1523 544
rect 1435 475 1523 498
rect 1721 559 1809 659
rect 1721 513 1734 559
rect 1780 513 1809 559
rect 1721 475 1809 513
rect 1909 641 2014 659
rect 1909 595 1938 641
rect 1984 595 2014 641
rect 1909 475 2014 595
rect 2114 559 2202 659
rect 2114 513 2143 559
rect 2189 513 2202 559
rect 2114 475 2202 513
rect 2314 563 2327 703
rect 2373 563 2407 703
rect 2314 472 2407 563
rect 2507 642 2611 716
rect 2507 502 2536 642
rect 2582 502 2611 642
rect 2507 472 2611 502
rect 2711 665 2815 716
rect 2711 619 2740 665
rect 2786 619 2815 665
rect 2711 472 2815 619
rect 2915 628 3019 716
rect 2915 488 2944 628
rect 2990 488 3019 628
rect 2915 472 3019 488
rect 3119 667 3223 716
rect 3119 621 3148 667
rect 3194 621 3223 667
rect 3119 472 3223 621
rect 3323 627 3427 716
rect 3323 487 3352 627
rect 3398 487 3427 627
rect 3323 472 3427 487
rect 3527 667 3615 716
rect 3527 621 3556 667
rect 3602 621 3615 667
rect 3527 472 3615 621
<< mvndiffc >>
rect 49 153 95 199
rect 273 153 319 199
rect 497 153 543 199
rect 721 153 767 199
rect 1224 169 1270 215
rect 1464 169 1510 215
rect 1740 106 1786 152
rect 1964 106 2010 152
rect 2188 106 2234 152
rect 2332 106 2378 152
rect 2740 104 2786 150
rect 2964 152 3010 198
rect 3188 104 3234 150
rect 3412 152 3458 198
rect 3636 104 3682 150
<< mvpdiffc >>
rect 69 507 115 647
rect 762 568 808 614
rect 1256 532 1302 578
rect 1464 498 1510 544
rect 1734 513 1780 559
rect 1938 595 1984 641
rect 2143 513 2189 559
rect 2327 563 2373 703
rect 2536 502 2582 642
rect 2740 619 2786 665
rect 2944 488 2990 628
rect 3148 621 3194 667
rect 3352 487 3398 627
rect 3556 621 3602 667
<< polysilicon >>
rect 887 720 1909 760
rect 144 660 244 704
rect 348 660 448 704
rect 588 660 688 704
rect 887 660 987 720
rect 1127 628 1227 672
rect 1335 628 1435 672
rect 1809 659 1909 720
rect 2407 716 2507 760
rect 2611 716 2711 760
rect 2815 716 2915 760
rect 3019 716 3119 760
rect 3223 716 3323 760
rect 3427 716 3527 760
rect 2014 659 2114 706
rect 144 415 244 475
rect 144 369 159 415
rect 205 369 244 415
rect 144 260 244 369
rect 124 216 244 260
rect 348 415 448 475
rect 348 369 385 415
rect 431 369 448 415
rect 588 447 688 507
rect 588 407 839 447
rect 348 260 448 369
rect 572 346 751 359
rect 572 300 692 346
rect 738 300 751 346
rect 572 287 751 300
rect 348 216 468 260
rect 572 216 692 287
rect 799 260 839 407
rect 887 420 987 507
rect 887 374 913 420
rect 959 374 987 420
rect 887 361 987 374
rect 1127 407 1227 475
rect 1127 361 1150 407
rect 1196 361 1227 407
rect 1127 348 1227 361
rect 1127 279 1179 348
rect 1335 314 1435 475
rect 1335 279 1355 314
rect 799 216 919 260
rect 1059 235 1179 279
rect 1315 268 1355 279
rect 1401 268 1435 314
rect 1315 235 1435 268
rect 1809 411 1909 475
rect 1809 365 1836 411
rect 1882 365 1909 411
rect 1809 286 1909 365
rect 1809 240 1836 286
rect 1882 240 1909 286
rect 1809 230 1909 240
rect 2014 353 2114 475
rect 2014 307 2044 353
rect 2090 307 2114 353
rect 2014 230 2114 307
rect 1815 214 1909 230
rect 2039 214 2114 230
rect 2407 303 2507 472
rect 2407 257 2431 303
rect 2477 261 2507 303
rect 2611 439 2711 472
rect 2611 393 2626 439
rect 2672 393 2711 439
rect 2611 261 2711 393
rect 2477 257 2527 261
rect 2407 217 2527 257
rect 2591 217 2711 261
rect 2815 415 2915 472
rect 2815 369 2843 415
rect 2889 394 2915 415
rect 3019 415 3119 472
rect 3019 394 3049 415
rect 2889 369 3049 394
rect 3095 394 3119 415
rect 3223 415 3323 472
rect 3223 394 3249 415
rect 3095 369 3249 394
rect 3295 394 3323 415
rect 3427 415 3527 472
rect 3427 394 3453 415
rect 3295 369 3453 394
rect 3499 394 3527 415
rect 3499 369 3607 394
rect 2815 348 3607 369
rect 2815 217 2935 348
rect 3039 217 3159 348
rect 3263 217 3383 348
rect 3487 217 3607 348
rect 1815 170 1935 214
rect 2039 170 2159 214
rect 124 92 244 137
rect 348 92 468 137
rect 572 92 692 137
rect 799 64 919 137
rect 1059 112 1179 156
rect 1315 112 1435 156
rect 1583 152 1655 165
rect 1583 106 1596 152
rect 1642 106 1655 152
rect 1583 64 1655 106
rect 799 24 1655 64
rect 1815 46 1935 91
rect 2039 46 2159 91
rect 2407 47 2527 91
rect 2591 47 2711 91
rect 2815 47 2935 91
rect 3039 47 3159 91
rect 3263 47 3383 91
rect 3487 47 3607 91
<< polycontact >>
rect 159 369 205 415
rect 385 369 431 415
rect 692 300 738 346
rect 913 374 959 420
rect 1150 361 1196 407
rect 1355 268 1401 314
rect 1836 365 1882 411
rect 1836 240 1882 286
rect 2044 307 2090 353
rect 2431 257 2477 303
rect 2626 393 2672 439
rect 2843 369 2889 415
rect 3049 369 3095 415
rect 3249 369 3295 415
rect 3453 369 3499 415
rect 1596 106 1642 152
<< metal1 >>
rect 0 724 3808 844
rect 69 647 115 724
rect 69 496 115 507
rect 466 430 542 654
rect 762 614 808 625
rect 762 512 808 568
rect 1256 578 1302 724
rect 1256 521 1302 532
rect 1464 632 1879 678
rect 1464 544 1510 632
rect 58 415 318 430
rect 58 369 159 415
rect 205 369 318 415
rect 58 354 318 369
rect 373 415 542 430
rect 373 369 385 415
rect 431 369 542 415
rect 373 354 542 369
rect 600 466 1087 512
rect 38 245 423 292
rect 38 199 106 245
rect 377 199 423 245
rect 600 199 646 466
rect 692 374 913 420
rect 959 374 987 420
rect 692 346 738 374
rect 692 289 738 300
rect 1041 315 1087 466
rect 1464 407 1510 498
rect 1729 559 1786 570
rect 1729 513 1734 559
rect 1780 513 1786 559
rect 1729 407 1786 513
rect 1833 538 1879 632
rect 1938 641 1984 724
rect 2327 703 2373 724
rect 1938 584 1984 595
rect 2040 632 2281 678
rect 2040 538 2086 632
rect 1833 491 2086 538
rect 2143 559 2189 570
rect 2143 445 2189 513
rect 1137 361 1150 407
rect 1196 361 1510 407
rect 1041 314 1416 315
rect 1041 268 1355 314
rect 1401 268 1416 314
rect 1464 215 1510 361
rect 38 153 49 199
rect 95 153 106 199
rect 262 153 273 199
rect 319 153 330 199
rect 377 153 497 199
rect 543 153 554 199
rect 600 153 721 199
rect 767 153 778 199
rect 1213 169 1224 215
rect 1270 169 1281 215
rect 262 60 330 153
rect 1213 60 1281 169
rect 1464 156 1510 169
rect 1583 361 1786 407
rect 1835 411 2189 445
rect 1835 365 1836 411
rect 1882 399 2189 411
rect 2235 445 2281 632
rect 2740 665 2786 724
rect 2327 552 2373 563
rect 2536 642 2582 653
rect 3148 667 3194 724
rect 2740 608 2786 619
rect 2940 628 2995 639
rect 2582 502 2786 537
rect 2536 491 2786 502
rect 2235 439 2683 445
rect 2235 399 2626 439
rect 1882 365 1883 399
rect 2615 393 2626 399
rect 2672 393 2683 439
rect 2740 419 2786 491
rect 2940 488 2944 628
rect 2990 542 2995 628
rect 3556 667 3602 724
rect 3148 608 3194 621
rect 3352 627 3398 639
rect 2990 488 3352 542
rect 2940 487 3352 488
rect 3556 609 3602 621
rect 3398 487 3678 542
rect 2940 466 3678 487
rect 2740 415 3514 419
rect 1583 152 1655 361
rect 1835 286 1883 365
rect 2740 369 2843 415
rect 2889 369 3049 415
rect 3095 369 3249 415
rect 3295 369 3453 415
rect 3499 369 3514 415
rect 2740 365 3514 369
rect 2021 307 2044 353
rect 2090 318 2213 353
rect 2090 307 2551 318
rect 2740 307 2786 365
rect 3602 307 3678 466
rect 1835 240 1836 286
rect 1882 261 1883 286
rect 2157 303 2551 307
rect 1882 240 2102 261
rect 2157 257 2431 303
rect 2477 257 2551 303
rect 2157 242 2551 257
rect 2621 253 2786 307
rect 2964 253 3678 307
rect 1835 215 2102 240
rect 1964 152 2010 169
rect 1583 106 1596 152
rect 1642 106 1740 152
rect 1786 106 1815 152
rect 2056 152 2102 215
rect 2621 152 2667 253
rect 2964 198 3010 253
rect 2056 106 2188 152
rect 2234 106 2247 152
rect 2319 106 2332 152
rect 2378 106 2667 152
rect 2740 150 2786 161
rect 1964 60 2010 106
rect 3412 198 3458 253
rect 2964 141 3010 152
rect 3188 150 3234 161
rect 2740 60 2786 104
rect 3412 141 3458 152
rect 3636 150 3682 161
rect 3188 60 3234 104
rect 3636 60 3682 104
rect 0 -60 3808 60
<< labels >>
flabel metal1 s 3352 542 3398 639 0 FreeSans 400 0 0 0 Q
port 4 nsew default output
flabel metal1 s 58 354 318 430 0 FreeSans 400 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 724 3808 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1213 199 1281 215 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2021 318 2213 353 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 466 430 542 654 0 FreeSans 400 0 0 0 E
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 2021 307 2551 318 1 CLK
port 1 nsew clock input
rlabel metal1 s 2157 242 2551 307 1 CLK
port 1 nsew clock input
rlabel metal1 s 373 354 542 430 1 E
port 2 nsew default input
rlabel metal1 s 2940 542 2995 639 1 Q
port 4 nsew default output
rlabel metal1 s 2940 466 3678 542 1 Q
port 4 nsew default output
rlabel metal1 s 3602 307 3678 466 1 Q
port 4 nsew default output
rlabel metal1 s 2964 253 3678 307 1 Q
port 4 nsew default output
rlabel metal1 s 3412 141 3458 253 1 Q
port 4 nsew default output
rlabel metal1 s 2964 141 3010 253 1 Q
port 4 nsew default output
rlabel metal1 s 3556 609 3602 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3148 609 3194 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 609 2786 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 609 2373 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 609 1984 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 609 1302 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 609 115 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3148 608 3194 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 608 2786 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 608 2373 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 608 1984 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 608 1302 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 608 115 609 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 584 2373 608 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 584 1984 608 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 584 1302 608 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 584 115 608 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 552 2373 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 552 1302 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 552 115 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 521 1302 552 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 521 115 552 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 521 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1213 169 1281 199 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 169 330 199 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1964 161 2010 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 161 1281 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 161 330 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3636 60 3682 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3188 60 3234 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2740 60 2786 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1964 60 2010 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string GDS_END 474074
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 465800
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
