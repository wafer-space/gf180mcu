magic
tech gf180mcuD
timestamp 1755724134
<< properties >>
string GDS_END 9502216
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 9253316
<< end >>
