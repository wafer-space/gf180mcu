magic
tech gf180mcuD
magscale 1 10
timestamp 1755724134
use nmos_5p04310590548761_128x8m81  nmos_5p04310590548761_128x8m81_0
timestamp 1755724134
transform 1 0 -31 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 359912
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 359598
<< end >>
